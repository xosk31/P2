XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��V��R+@���Lq�����*��}����J:����C���C�X�N��"(,+��TR-�}�ۓ,7<�	(C��UG��~��m��"�1�f��?�B�;���x�~���?k���ha����j�a0�h�|!Nn���a�J��}�V-��� l���y�ß��q>���,��g���.�ɶ�9ç��0�<�DS�$6�����[��-+���"FK��P�y���,]K�wK"�#도E�?��� �\/5<�dU�t��)����3A�m.��	^lŉrn>����^���0yl%W}������b���b�N]�t>|��Ht���x�opB�͠_����t舦���n�6��C���L���
J�Z�\��J�C�R�xU`Q��'� }�s���� 5`��5�PW��Y�i��-��Sz�8���?6:�wf�c��
��0��Aw�]�]ٙUPm�Z.ۆ�}"۳C�H��@����$��4�nxuQe7��d�;��{%Ĳ��7A��D������h���p,S�}�ch��3��x��ա�[��H�>���>iI�V���<u:rI©ܩ����~�_}�	��T�$�����Aa������&���۴��k�cOy,�\�؄&�/��ɋ��Q���z�2ϯ*��p��X�vg,>D�h6�t�w[m�WV�_B��&=�|��M������n �sFm���?�H�2����k��xf���Y�o墒|CQN�񏫵�Z��XlxVHYEB    29da     af0��	����J�=f�T�&�Q�M�DO�+���l6�N���(��Јx�mu��t��_Ӈ�\�u��D?rV���
��ܨP�bqe�Y˶o�g ӛ�-K�O��(�法�'�Z�t�**�f�b�t@�E��?��>�i�~C��r#��ް�W��̓L�# �KZs��[��e5�c��>Rz���c���]����l���L[��K��tg��	�%9��]�7f��N���:!c�ؘ���E���<\u��T�D���5��|(�׸�̻��M���#�hW<GkbH�� S�3�9�n�!j�;T��o^Z�AJ�a�"�I�:�V��#� �Cc��,�I�����-��U�.�\�Po߸� �^�5�m�W%w���*��P��ZL��h�x;���-��3,L7�(��4�D�%�
���E���p��K�ss��:���-��!�u�S�C����uȴ*1T'w�v�Tm�B��Wcu|m�k􁸗�#�^���d#HQG���;)�p��t�'y^=u��isZ�1��*�,���Kýj'���اH伈L�^d����aW9���
4�ʮ9{@������Fu�/�.yI�]�N�*z��+Ao�e=���B���R)��pQW�� 2��,�O���i�n�[����o?Y�G���7м���C��Ğ����#�v`�$�i"V����(�.�ޖ�@
��xj}�`O��sJ��>.9�M�NB��"�:�N���ôE�F�")+��U�=�c5mt'�|�W���o���e2+<���#k���v.Md�a�:�J �^3iv
��rO1׭�e�[��
�B���_�6'gw���w8h!.������W�S� CY�{��r^R(Sr�0^:R�(����\Dz�~8�a Zz���%9��k։���=��%0p��F��z0�7�:Ga5��7r|}uԌ��
��&��
H�[�O�����NG=۸�	����\��;sg1}�w��`̯��?���ȉ���_����n��������|�c��ۅ��,��_A�&��Ď
<Vu����-ҋ��%�}+��\Z3���h�[�}��A��C�nQPh�ΝK@(#���5�B�8�8�Z��7��u��ŕuW����pW�)k���
���&S١ʛ3tψ��;��#�4K:e��U��g���S�ö��-��Z�ٷ�Dn����V�8��%�Å�HS�FL_yT��͉��<[�����L���#��L��ݵ��m���!�0�8���D�S�H�1z�rg�^w<�s��b��������>�n��qg%�0T��������E4o��r�4��r��k��)/�@?�p�E/���|U�2p��VF�Q�dz�z����u#M$����+ꦘ[qD�|�E�	���J����V��K��Nw��.��h��K��o��R�5@箰�.���nbQ�xWo�C�u�=s�xȡE�B
^�Q���xA��� �p#��S��8�oм�Y
�cw�Ŭ��n����2y9�ΗT�gѴ򥉇�8� ��V��l�,M��6e�Cr�aF�Q.��|q�_��AZ�̝O�j�l�7ù7�I�� s�V�J!B}�3M�hq�ف��`�&*NhRꩂ�
-^u�������(_���qʌXhnp[�1�n�\��P�&�����m�Uۖ��	�6�Ek8KuZ(�`����<<=.��ۃ��g )p4g�	���I�uv�a1�nw"e���&(!�#�`�,� �u홾�y�'��Gp Zv�/B��fX2���.%�L��`&�{W%����V(e;�c�������9�/E
I���{�C�F��)T�zH��,�چ��J��e��E�IҠ��Q��PKa� o�p�d��(m������ş�(s�uL���V�5��u�:(LF�/ F��O凉9��`�c���t����T5^.���P5G�V�hf��d�n��[�*�c
��w8%[�(-�E *ȉyRf��Qe�x���t��+|����3���TG(����[9 �>��dgi$.mk�hp���2����(��Xe�B
���� �����w*�Q��n^+�� �~Y)e�dcH�xPF}XA��?s=tfz|ւ� �X�Ƞ��zG݌S=��]�!���{Qr�N�o?'�;���J��&�e�>#/�����u�z5t;��5��(̵,�eK^�����(I|��F��O-ФK`����;�Lm�}��C0�d޺��s�Yԍ��6i�YOJ��7�\?K���N�*��ᛘ p��/&Ku'w�՘G=����-���C��O\N�)h ���;��q�Y��Z��ẉ�JaS����g !��`� )@�,��ϛY�"*s��\���SXW�Hl&��>5ր�ݧ�&Q3� O/���"Y��3�Y*���7V�D��r�{���NAb
MO7���	4����e=T��!23������-Zۖ��kPKV�4y8�f���o^��U[����ʧ�Z��ĥ*�h�Jv�2��Ĺ��v�a7ѶL�;�]_��V�ᜓו�;�A����dL ���H}�̈́��tQ6��l��'�N��`��7i?���ѐ��0U�-o�e�\��w:�)��؍?� ��4�^���2Ic�uG�p���1�0=>?o��`;EuY��T�GG�����C��ԟץ��Q�*w~_�W}�����p\B��i�������"�6���,��<�6