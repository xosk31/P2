XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��N��b|�ay�}�M�O4ۿ�]�'�bB� AP���ΐʤ�e"�����EM��ᬥ�ŕV��o��Z'�z��F�eӪ� ���J�RH�[N;aSr�/�@�W��{���R�"�-=n�&y2��<���	ׂ�	��ƒ���E6ޝ<��F��P�;@�|��?�yU<�(
�C�J��h��X�w��.��c�ۨ�* K��B-�io˪��Jk�p!<�3�ș�YBǔx5՛Ù��0=���s<�"�sR����'oX�����}��{����*���#����E�ܵ�1�����$<��"6����#eېT=�<�D�(�}����ZN+�k�ܳ������B[�r�em9[<轛��h��Ā2�����Ax_��ӝ�{�.�3�,��xӛ�
���TG�aH*�k?�fKq��kTi�֔�'P�s�8�,)Q��|19x����<]6���e�t�gh����~i#�@�_?I'��Dk<Ʊ�P"E���buU 4qP����E�PX��8�Q$��R�h�����M d(���g��ҤtG�	M;� %�.TƼm��ķ�W]����ۗ� 饻!l�\
���4|�ƵV�i��U��*��._t^�+	3�@O����W�ݬ��bNx����XU�"W�K^�j>��H�^t �?��]�]������� M�s�����z��U[�Tҋ�҄r�.f��D�CҨ��
�|�=��o��ɣ�-q �E6�[�K����XlxVHYEB    37dc     af0�/���	��C��E��U1��G���=?e��X�-�8'&‭J�H*8��2��(����A�>�J��� � D<#�L盦�	w/80�z>�}e�g�d5.髊�%b�����խBf��(zI:�����e������{���|��)IZ-��zQ.� _�*-����5ox��XNάZ�3�/��Y�n��!���  wđ��0ԋm���S�����x|q��`�4���A��ѽM��Z�S�Q���1fΏj��.�T�	7��ʮ`cP��0��e�jC�R�-��J��	���uWd� �ֈ�62���A# &�DK[�����
������xݚ�R���H�)��BgK�T��)�kh[�ai�P0�����p��y`0�˼�fK�qqw��۷�K�ɍ�
��*s%�7y��R]�����6�ayڶ�z�E_�:�G�V � �5vViz�?�����hAd96P$\u؅��kH����UǞ��m�9Q&�a�>�C<]�
Y鑐�	q�w`��Q����,TR��6{+̃�A�[zPP.�oٗ��w�}%��^\"�E����P�U����fl���U@YW�^g�S7���2�<�D��D�kU�r��������?L,$��L���M��_�������7N��EAc%���5������/EH2�������|91+_)���_:�M;Ge�"����b9��'�L[ಃ��Q�ȵ6�U�77p�.>h5�u��,&D���������h��_����Zl��ɉ��\�%��!M��'6f�Z;�i�ƆI�&P~��U�ؔ�On�B_Ό۪k�Q^����=$AW�"�n���Q��؛�7�9��	~�k�/��ٓ2r1��/����IB��˴#{"3�'Ա�JԵv�Ik<�+�G� x��Ӟk�1W�*��֒g���B_-/�ٸ���|�ך����F�Rs���/���b���`�<�5�t�*Z�z]~��z^8ͤ8���񏟑�'8��;����k��c�.�W��-!�V$='\��"?��B~� �mA�KD�0�|�7���u.�����m|Ձ�۝"���MX�+�8x4��8Oz%XF[�U�����ʒ������K��_�����o����)�#�rتqz�#dXMH'V����	�Y����v��d#���N��~5O:$��=�ȐȐ	�(�1Q�b�*<F鼉>���5�f'{�p�x����d,\{���*Eҝ ����?x͐�٧̍��׏փ��<#-6�[�_�ɮ	��tt�ʋW�L��W�Nj�{4�C0a��aL�7S�OҼmX�Kʢ���r(�йZ�����:C���Z�኎ˢ���� N�>�a�c��-Q��y)�k-Zj�/e�n�e���F�{���+0��M�N���D��K�a�w��LƱ�մ�j1}-��Tg_�Y����o�Ck�tɜ����(ј�ɇo�zb,fc;ӽ�铞�Ȅ���G#OAD0����5&A�k�zKҋ\`��zw��;z��II�	<!'{a��;�*q�_��1�{g7�iH<6G{�&�f֌l��-+	�X�>�2pY�*N��f�*b�}z`Dss6u�%�� :������>(�^
W��̱�r�o-y[+n��NqQ�v֭����R�ULFʍ���;3 �.L���f��ML.�~���Ѵ��"4�ğ�/e�p�퐮U����CU�4@���}�3D���cՔ����3kjb�x�����-��ս��[vb��j6&t�'��dY��-�������C~��̾	�'�$��&u��!���$]��fy�tɷ��;o�e/<�
��	%�E�?�#s	N��l�.�i�t|�^c�/��˶W�d(�������G�[�d��f��mr4)hk��g����c£�h�����~�~	�8r����h��bz�S�0Gӱ��^�>�I8xB�[u��5e��¹�������G�(��=����*p:Z����k7U#ƕ=9��_�(��ÁAì��DQ��s��\�a)�������\�{L �8yj�(	���`���tf
5z��V��ǧ��/e�Ž�F�2�����S��>2;4���y.|��׽�V�9��&(=Wv�j��OqU@���U���x�-~����<%�d�K�4~�{ jk6��z��MAF"�eڛ�.Ç���H�ߨ�p_�.i�.��o&KR>�Z�0᪕b�щ���ɡ;/�Iu�)�̱��x�G��n�A����R�:!_`Pw�|�q�E��3c�nmc\�`��Ő���SB�T�O�o�"7���k�I�(	㱥
�?���~gw컋�%���c�̰�|I3o�#xУCLȱ�4��sw'w�m�n�+0FB�g�ݢ�=p�G�*޶�Ut»Kl,����z�+��T�˱3^a���Nk��$)�C��ɮ��g����׉q�x��x����P�O���@��l�*)�ɔg�C:�&��c�9ƒ��|�Z�Az��N{�.���A��_�=��#E��)�wj����ۑ0k߭�R O<^l��+�;��6�Ӵ`�i�p��%�g%��
�Z����
�Z�R�'}���gv7�Y������9���6������p��M��J�	,�qB��N@l��x���#w����rT��,hԖ�r_3��� �~(g���4%����
�]�d���+�}����L���H��(3V�Oڹ�b�2?