XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��$˾��vUՃ�"�f·%R2���˙ژ�|;꒎y�u�'f}l��G�B(�FN�8*�}���Sd5���
��;(��+J�@0Em�${�F��
���Q�
W���s�4�鈂��"�v��o�<�.�d�ߌc�/{��x��-�px�~'o�a�C�گ��pݰ	��9�9�����u;Ţ�E��%���{>юs��� �!��Y�Ja[C��fA�٢59ξ�8RSv5�I}�Z���q)L�l���xU[$J8��]����!��>_����pR5;�����X�wm3w9�x�R��KL��ϡ��]�
���#��%]런�m���0\��2�9�bv�h�2�kN�|?�9�,������?�fF��=�U_�a�_��4X���	lZ����<<�F9�dp��[��6�&j �q�f�f�D"�B��%�V�ya�b���jJ]�
��w�(����$me����'�w��%�RV����)�A/��@�����|�� F�Zu�>���M�I/��#��=�z��?C
 �ߨ�����S��$
������1�aa�|�{��SԺj�_d]�8�t�=��/���Tv���	�$V�	�e�l���h$(R�"W�SJ�,��A$mm{0e3��N()#������m��谟5zNP~�]p�������y��`���&�F������a��g�N���{oT��/
p��������(�L"�_��?U�^�\��m�ۛV*�zYhDlwm�.��[V�<9.ZlnFE�G�\�a�:XlxVHYEB    3504     cb0/YJ�E~�]=�4�>�0@S�.�7�,C��J�vP~OwuDj��I�Q�,zt������ޘ_<�tuY�m��M��jq~�����ޒz�"��`�,^�S�2�.��@��H|�-Tl`zO�shrޫ�%��/w(:#���+�"��L���U%qAt���m�n�d�ǜ�9���W�-a���U���jR)�GY���=|�?��U>�*a��(+�������t�wlM˕S̋��f�X��j��]׬��`X��)Ƈ����ȯ�W�!�Xb�f@U{r˼�<��a3�ߏ�#��Pb���i�yr�|�4��=c���
��9Y?� *C�T7E�6p�n��Xn� �~;�`����.c�S�����ĺ�F��[�1#:ڏ�����+n���/=*�U-ل}%_�����l-��c�?����Mc�n�߲�_lu,�ϋ�n�Y!fMlL�\X��.J�����f�Us�rW��×uD�\��;�����3���4*Td����J��x9���R�I���t�6����}���.#Vj:�X%;2f�k�qp7�l��I�~�*���6<0��Z_Or l@w�D(Qw��%�9"f��z)�r���Y���jU����K -�}:I2�]dûMV�L.�q����lX��=����y_�^�m��c�n.�����.��r���U�]�23
�*��
���.-jC=�U՟���ݪgy_f�'�W"��G*�Ԛ�a
8�BqR������Z�(W��E��I|0=�r�v ֬�Fp�Ő�*YJ��M[C��y˚��G\s����T�r�����iF��'/�*��f���0��ϸ
�m����4~_��D/�-*V������F�f�"�Lb����ULN6c��I|�������H/�t����͔��Wu�(fkzx�k�_��9U�ȭ`��8f8݅f�X��X�+<��I�J�
�x��{E�T{��4�E��I�xn�;��H��x�ר�i�s{7��o?vM��&4B��^��tz��R0J{�z�����ԦB�/��l0"!2s���ɕg�t�~��~z�5���F|Q;�/�9|��x�t���F��谬�IG-([�}���[l偉׃���Z�S�ۮ�͊�\�E5�"7�6m)z����yUFV�W��pΚe��.�K�\#V�g^�%���)�xA�p�G���Ĵ�bw�1�67ڈ9�sh;-�0�ף�|o�È���2�ڪ�P� ����O�vUÐEѡ�3qV�������y�b�b����Vb�Y6��1	s�ª$C-g��;sGwƲgs˚[�F~�Z"�E����A^��
k��*sD xo�C<,ͭ�^@�P�l"��o|�u(����{����,��^�ϐa��bƓ��&��|����h���4�S�0E���oY
�`46z̩�w��_C�Q~ s"~��ʼ��Lu6�����������@fԲe#�̒ғ������B͒^�G@�D9z�~�p {�!�Z��:�]�K��
D"m�C1�:!��J�s�*]g]7�e�/��Z��β���b<0�I9��ڪ�jQ����@��BʷN�:��~��.��j��]��B>1�a��翀�vv֪&_����D%=�۾.(G�"�CS
%S���D�g�A_�I]����9�f��\�tC����9��L�Z��@;�}SZ�����G��n-���wG��m?\5#>�{�OuK�bg��+����3����Y�(�?�~.� /���j�����Oѓ���\���e��!�2#�O3��O����8R�L�r�і�¡� ���r�t��̓��8\�J�D�X�I���企8(䘤��Wο��������\�h�����V��,��;�A��s�����-N�7z2��/�������^ŁUL&s ��A¶��' �B���Ks�b���$�Ӻ��c��E�J�37���̇�o�=t8��РB�����y��^"v�Y[�\ζ��GG�.Ka�b��b�A����y��2j�W��$AV��f�e�D��-�$��sD�����[�1�I�ߨ��؇>T9Wj$�'ͪm�V��}�@�I�<!����f_^����L�Z�ݶ?u`���Zv�f-o��5e�;���s�������W��k���8<_w�g-t>���U�ǨRtF�c���)�&4P�eFn�KK����(��ǽ�aԏ5�5.{*l����p�8�0��
T;rE��@���zZ��g���X~�Ed�/�M��y�i�]�&�s�$�R�!c��ꃣ��Q�\�E9�7�[$�-a�L�.��N�ψ�K7yP���������ŗ�)r��PzK�H8��������%�-��|cp��Ӄ�`7y�j)���
����9ӫJ,9o�*�1o�4��R}�� ���*PP<5E���Q�g֛ȻɳR��tb�b�ϼG��R;l@��� Y)]`���P�U>��v���Q���cl��)T���%�v��k��Jq����HK�A���zh��j=���F�R��Iݳ�FC�0�Ai��-������{���ӹ�|R�U�5[�5>C/߭�M��j)J�K�\�M�+,~LF1U��Mr7k�����o���k\��� �đOq�S��	��z�Q��I��Ȫ��8
�+�	��6���\�O�˼���+r� X�����˒�afd�H�F��{�.q���Hn��񙚠0�9ߦXrGU���?����!³�$����۱��f�U�U?(dn{�d�D�m��?���%��R��M����e��m�v3�5���d�{��C����}H`�T~�1R�0*.�An5o2}��6c4�'�y�)�c�������>'qf��va�#�ۜY="�n�9��5# ���\3�~t��s�y|s���$Ǥք��Ҟt��
 o���ޟ���;d��P\@}:�>�ר*��Xbd�Lz�)�a-��L��}\�l �e��n��P�¡u�ۤ�pӀӈ�Ĭt����޻FRF���-��Ѷ��`��Ħ�)�۴c��Y�5�%���=~7����xV���-���n���_���$JP
|��d�yd��z�O�|y(xU�=]�Y�;���1[`�N���RS7H�\���E���\�@q��jB�ae�Wgx�N�>����)ExbQ�
�E��Z3��0vD9�9��?g1z1N�