XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��X0bp�Ǎ����GAR����6���l���I���rL�xeu>H���;w����A�=c���)��d��b����*n$��Qb���+МH�^Cj
LPi�~�����7���HQ��q�x�_�U�|��*\����V_� ����h]+�2-��	�@1�% ��{aBZ;�9x��aa���8�����w�kMY*޷�@gR����GJ�9�0�N*o>4;]��8&Ҝ�̡�ht˱�=h�&S�R�b�pM��<z��;r4�K3�\qz�d*��՟��8�Uy�,�,���Fj5���')�0_J!㾘M���HGQR��_+S�kN[�4�o�P�c�r�.���6#H���i�{���o��gD��/VEj ���}�u573GlMUY.OI�����ED��߲;�o)��>y��(ik#tG��V�+���GT�z~\6��=�����S�ߗ�:����T-��ag����Vj���O�a�~���`�%S���=�b�@Wʥ�R�>��
N������c(�B�6Z��ho)T�'ϖD؂�6���lhY�"�_F���u�g�:l"���pRǴ�o�r���W��1	�Ep�6#������S�q���=8�P6.���CJD�5�ЍP�!_:V`��I���S��=����s�;p��(*�FO����P����ߒ��fa�����m���B�2��0�D�\A�61<>�x�ܥ�Q�Tmv�S̰�M{y�C��>�Q�XlxVHYEB    fa00    1ca0��u�mH�f^�kN'�Ϝ�]�^R0b�2i�/�I®�.���L�S:SZ���m ��z�8��%��M����Sv���9X�7`sS�:g1
�a1j�7�]�:�c�R�I�0��(��F�`�|b��C��[c;�>�G�p��~��<�LH隽����nI��/��-��ϯ���ēK&<qE�i�M���f5���XG??y��J\���uS�-E�;%\����r�k9�]F��=^�����Ĥ��1�ږ#WG� �v��50��)\�'Mk��O��}ϫr��7�)H����ˉw;4ݣ��p96�R�R�P	ܡ-U���ޞ�P��Ү�x7r}��S�ݣ懺8Q+��o��KTN�g�y��'N��}��YSkEG�l�����s�g�J�H��{|�fY�?��������3���m=w���W���]�:�×%*67�Ô��1Lݷ�����ʦ�g7e Q |�\��1�T��f�_�|"那/P��qܘ���̄b��z�+����?�Z'��}��q ��&�/�6����+�cW��z���[�:��Rt���u��eI;1�R� �n��c�W9/��2�a	�%��͐PF0l��]}�n�,�3^�g���z-���pƼ�]�g@�Lo�p��r�ͭ��㧱�t���J�5���
�B��g�ۊ�˾"��t�fc{�E��Ѱ�Bw8׵��S�޴F$�7U*�G�(�JbY���#����H�<�ֹ5��jX)������;��l#�b��F� ��0�ϔKQ�:<�4��T��|��Tm�)D��`V�-d��Wo��G�����T"[X�ZD������f�ۨ���I�bZ %�.������n��������jR_ti�zQ���9��\�Ĭ�<q��٤����t y�y��m:�r����ڋa�ޮ�N��p��
�CX1��Sz2U�S�(7��Ex<K�pSof�j���`�5���ܙ����7�nq��"Ɗ>
_/-[�M�$>�Z0y��dX�/d  0Yc!W���q����"����+<8�d��R~ȏ�h3+��>ȿ�_Ls����m,9��&J�;�˺��,o�;��<����V�Pm�nZ9�K'��N`m� ���˦7�O�:�\�9-�X��	�(ؒ+�Z���� �[���oeҿzYma�rߨj*N �BU�|T ��݃��@U��
��V_һ�F�I��Wqk~� �N����P�k%��QO�A�.��]ѱ�ΔF1��h�	@�>HO���ѡ�a�:K��1[)N���"������R�H
����J�
�=�����,�E�T v��H6<bBƬ<�C�������E%Yi�~���@X��rl��!$":�l����� vZ��m����Z�4�b�/5ݫ��ɯK_-�$��gi���W�-C9��q��VW�v�r-��⇀����^���b��4��N��K�B7���5�e�გ:l�T$Eu�/������������8��6�qr��ʸ�I ��������.���-�'�&?�~A��$��6Ǯ���υ��<Gg蕥3�y�:[�����H"���F�F�ͯ�Ĉ�p�Tש�"�i=*n�ߖƴ5E��E��@�o},S_�| kMa�X�|Ѥe�W'�'��"��u	�6+�"���'հn�eV4Q�	�q�>��RI��� `cCu�'�0"�7w�{��+���9���f���ƣ�">o�y��H��`�^������l�5�2J�o^�3ғ4Q�ͫ���v|��N�բ/���˷C/536�S�H���K��c����y�k�������d�?F�	�ޥ�����ϟ�7n������+���7����<5��Z�2�����-$�A�H��ٯ�i��A���%A�$�*�@��xZŅ���:�!��?�h��(1� ��Hl��+6�9/�CP/��Hl����Xpv�Oɣ/�xQ���/�L`���Ԣ�ZJ�E�%�G���v%O�6�}sKt}!Ao~�踏���VOb֖�<���F��4M�c�'���H~R�	Wskl��@��w5�k�i*������%S�Q�}fj�_�l����>�� & ^�%(�ŧ�;{���I��90���7N��S	�\�0�ء1\6kd� 9��a�-�e��<87K@Sb�:Ѯ=�Ni�d`�ҊuM�*?������3�!G�/�d� �sǵ�J�?U��/1��ޝYyJ2j�?y�PА���06�8���HqbhK�{���I�m��rt'��{�u������) e@�bOT9afKSD�V�yr�`�c�`�KUڷ����&q���ܵS���X4�lC�ː𼄦&�wyj��������O�	w���}/S�8e<&����#��o��������#�5s�E�=8�(�9k� �-�0H=3�, ]M�<�-J|�ѧ�+���MuL���?D�a�l%̥�"{�S�x�*�@ �%@lA^ڇ��T����5�5�_ =@�EΞjL�G��@FZqQ�E�wM���t�#��S��2�|"��j[��F���G4m�_�#-���Q��ޡ;�nF�?��M�L��]%m?lg�����{.t��7��թ�:л�n4��<I�d��n�ɕ��f��!�"�e�Ӣf�����χeΟҲ. ��Pk��(��C*!�7�~�Ӫ�U=�[��C}S����T36��ڎ���2]+�(��uR�O�%}C��HrV~]����/��7?���m"4'��p|<&�ɑ�,⫀ڔ��ҩlZX���n�[&a��|��.ą�I��prw��5}���Z�XNM��9^X}`��
]�ٍ�!���u���+ 12~BW�X�E�*�����3��_���=6�&�B��PS��Ȑ��w������J�)����<�*yw2+ �y̦g�)pC^����KG��>Kd�Rl���}�m'p��w��:O
�)��5�t��?�0��zɼ��E���yQ���E�G�\� t�oZX�ymi%h>�3��'���{ֿ{t��Ī9����
Jؾ%GTiE����'�ۺ\�qH#���Vd�Fc��-u����[�P`S�V�խ�;"�-%·�9#��z�^&�N���DI�(z�A��r���ݪ���z
#5?��,%������/ ��f��>T@婣���A��r�M�5�r�lr\b:��w���2�e�*x�+�0�k^w���_Ļ�	\q�a�k�\?b���Pt3L��G���? �=T~�$j�����LJ�0f���Q�6��'�^��t��p֋�9�ɾ3%�]𷐞�/���`��\�YH��:d^>����ЉMFV��B+车�,)�$�o��=T|�)�����]�1 R
�=��u�b����S�Km����C"�[�w:vz�A'nk_ܫ�"�~�QeEk@�|(m!��X���t�F�~��J=�9\b�}�/}a�'�W����(���'��}��zO^�y6��!�٠P���l3Շ�`��^���[u��D��-:s��(j�����q��>�ؚ3��K�- 2;�C�Z���|j� ���B��b�)vo��%�J�i���Q�k�.�5�H��3C �=�d6���x���V�t;�C1V@А�<x����}�T5��b�b����e�*G��Q��!�� ϐgӐ��-'������VtQ`ˀi��|�%B��7s׌��|��	��c^��M�mER:W�Iv�gj���v����ѯ#�����x��=_�ŏq��zm�H�hS�'��j�֊�Ǔ��N6E���1�n��9�N��R��F�8p�d��=BW�B/���F�k^,U�@�n�EkV ~�RR��޻����y��A�.V�U�h����Q�قn�`B�A=8V�2��M�o Dٱv�@�^�~j���7P��f��
V ���b�y/N�a#��H2L�V�▦��oZ\��/����|(t�����gW���ث�������܊����&��6 ��8�!
"�[X��]�e�iq�l)=����6��w���W ʵM��E��}�w�sIR"Ɛ��G�ډ�+}%�0I&�v��O"�ĩ���k\I�at���·YF	�җMh�S���A���FF�io�ޖ@G��-��+����2@��I^7�Q�a,׈w���E�/5������x���ï�ktВ��$XĸA��DY���X�o����|��e�v�������ֈʀ�-�HsC��#9��̰5G�v���%J�ߠ{�ψgv����4-Q������&���%��0e�������V6��qՍ��T冰��b������&�V+��e�v�	�u�/^'�x�x�����`o^@�	��b�zZ�!���L����u�t��'�
������o�DN�Wf�G�|8����_���C��m�c�L��n܌���_
N���Rќ�u�(4���wV)0�"![�sV"c:Ϝ����bnf��kqj�E�)��ʼ/B�����|�qSfߩ�k�&:�͸���k�ʋR���caZdk_{�B9��F3P{����;�t�].����)��fV�be\�Пk ����A�����|&��r/���#�RŔ �[N%��)�q��n?�����U?n�߬V,M��x�<3�j�"=��D!\��dt��&�o���E����M�\�7����.Dy �J��X��ɹ����#�C�8�e;�V��:�(D+�Sǔ �2���{˿҉Bާm��Hm�!�:l�*Cf\dg+ݿN|���%��U��]�$�Z@疢I?e?�%�ӪH��c����%����V,G����u=���Ȥ���X����٣,��lЌ'|""�L���xA4�j@WL��u�]�Oi4���ЭM�`c��_]p��Dѫ JB���M�I�J�bVVo��`�Exw��r�dya���Iˍ�$Z�C���Bsc��մ���c�{��+�sz���������>�Z4����Ɓ	#%6Y�M���	�D��R��/W��Vn!�W���ִ�Hg��C�1�G�"�\/�@��;��־�T��C��(1�k H��V\��\��S������$�Q^���i�U�	ī{0;��LC�u������vuRoG�c�k������t�.����m�&=�>Lb�򎽡�n���@�xj��F4����y���d�� *�F�u5���pG�T�5=p"�SL�-ι���群��N��n�^]��4��c�^b���N�kE�rswz�I�/t��FѢ�F-�����y�����In�G#O]s���7��61�=L���ȮHeZ������=�@C�_
��=�S �;	��,��W��}$��fI붝�%B&J��V~��l���6�b�hj:�{)�cX=�#%�X{1/�mH�;�s���Øg��BWQ��f.ܟ ��k�7��J��bnI��=��dI�iV(��|�����|/���0��r{�u���AE�KW�Ͱ��89>1��h���.���Za�Ό[���&��M�P`�9� ��ؖ��v�t(�x	AI��1�m ��Ԭ���3�u:��Z ���^,ĳc�,�e8��,�,�1�)�?�+�ׇ��~�,�-	ϯBA2\}o�����d�@%�ջG�N˩$i�������m\�a ���N`�
���sp��aH �	�֧�~� ��^����ʏX=�#�q�q��[���@��7?K��a��N��_{�~�M?g��>�Y~w0APz�/<�v�{dI;��.�{��A��9w�n��B!��y�-!��䒈<~����-^�`r�H~��k|���΅ �8@���S�ym3K��8�Z�/m����^�j��yQc�_��y�}�~�}�o�>��Ɲ�7-�y�¥a��Z��]�`D+��d`��0���`�"ݙ�Vd�6А�8KEw��E+47��@ET�q-d9��?��r7 P3��>n�P��M��r4\���ꀢ<{h�H�f]Ѩ��?�)��1�����q�=w6�v]�WV+U}X�z��js?��cd[o��:��8��.���V��Y(�˽���١�d�mO$�$��3�2��נ�L�����6$��hg���U�:�n��k\Iw��e����A���
̅uk�F�c�$����EC�����/:�LI玤E�l�*��s����nBj���#Gxχ�Ig��XDg�%_�)'Y�e��>��k8�P���Lj�[�|�P�`T��y$]����Z\	c�W	
��_{]'�� ��v[��ZZ�E����ZlH_8{{�{�Z�(�%'���v�4v��".Z��)��)Pݓ���d�4֐�� �2n`r��G#�˜m3^mk2��?���ߵl�X�R"�+��C0�K���Cf����u�������.��q>�OUO�x����hO���_ɕE��>Ʒ�RI�\���Fvv�ss����m�a]�;�{���~bi�b)�n���T�p����`��=��Z���ڪ�1�w�zl)P��!Y��[��v���r��;H���A�ځ�l�������$:�>#�M���"(F �>�H�u��L�s"3�&'� �rs���-$����[cm�T4;po��R����i��2NCy�'v�_~!�ؚ� ���ОQ��fq���<�mx�WcVz���QnA/�t8_&Nt�Ψ����qٙD�/f�lCHO=�p�ӧ<�RuS����:v����S2%�BB�W�6���F%@�����W�:f�4���Lz��`0�E��tS��\^�Ib�.Z`cD'���:(>��h\��-�1�SO��%��'���_C��Gd��B"��}�5�m�# g�b?a����p�Mƪ}V�qۑ(~�ڥutn4���t�6!�r��((���[��<,�t��}�^O^�*¤�JU�ݞ=�&'`���@��K����MY�;��uSɹ����ej
\����o��`�P����1��D�ü���0:DF��)�_�ݟ�p �:ڋ��S�`y��v�c�C�+��:ѓ��\.w'nQ�-�;~]Bm�I�;��'VO|S�ԟ�W�H�JV]���
���4��m]X/��,�>"����{�A��$krP��>���B(�-Өe��x�`�"���Γ4
u"F"���`|��iEXlxVHYEB    fa00     cf0��*6j�+�`n�,��H~g�uLC��Ƒ�Q�B¡xt�3	�7��+ωؐנ���~��mm֟�yI�"ׂ�T�iF�32>Q��-[�zr�3�����8`Ol��pp�+����|}`��{t���U7��&��pa)t$���JÆK������q>64c���*��*G��W6ë��ۀ=MR���Z��79�V���CN|���M�	��jiظ*�#U���l���(��>����E��F���W!�f��D��0ė-3��6×:rcZʻ�(�)�68���WR�ی]経|���m�ug\�p�Β�ܞ �pU���������!\��DBܵk��<������K��[�.�,2���f$��}`��?��U��[(�AľϪ��\:�Zo�Π8�J�4;g+�_�{�h������+�:�0PR0l��k�<w7�7�~ �gª5E
/�UK��d���m��n���=Ơ�'8�J[p�ӭ�j�4%�[�X
�0�<�@؇�.5��f
�e�%L�/y�)���p����!+�&�0�zX�'�៼�g�L�}G��v~/П�m\3�,�3���Sk��Ӯ���3a=��ݛ�A��Br>���w�(��7c+/����)�8���-�h��ݷpK}�6�����dW9þ�9L0cD�Yw4q��bC���>QxW���Cզ��Ƞ�f~�H�E�������
l�2�k�����Ӽ���������/f��!��j��'WSw,u�S�a,dbG@wa.2;KRY[a4qg�=y,f;A��Uu��3����qp�"o�4��\�E�q�ڼ���֮ckc5"���t$�= co
*���k��.��vTA.�	�-֌�Kz%}m����*qfn��� �.���9�]�]���[�����2�ӭ_4Mw���-�/�ŸT{�%[!ؒ�}ɶog��/�N&��U���:��	�A�6��#����I}�l�K�}��,��6�5�����G���a�-��L���%�����k�]��Jh��o�gSAZHdD��.��_������x�F1�^IM L��U]�RQ�|@>CP�4�y���g�q���ƽ?a�TA`�ߑ�B�`�V%=_�KG�o�w��I���_S�@Dl�"����Zce'��'��S��8w)��&���ʳH*�^��C%Dg�<wMd#Y�n�?-r�0�{��_"�U�Yq�A��a�
b�:v"}b��r `@��C���=x��$�Ft�f�^�j�T���7�bz�e�q˹�B4^�����ȶ}�'uP�I<.��x�4�fj�HS�c��w#�2�=�S����+�-E��V����u�_ʗ��:n�{j~��?�y3#����l���p�N�f���u���&]$B��"�Z���֤��A��d1Wh#��3�1DNc�ݓ������<�A��'�W�M�/c�;pw��Gi��k��)���(���o���H#GM1D�W'���1�͍n������T�'3j�5��0�U����P����7c�DM� ��K)��H`���ݟ��������s7���2z���~�D�ޘX�x���x}�U�:���фT��	]�� �� �UӖ�$�nq���%G%���4�p�$zw���z�lR�a�;�fҪƂ����6Pv�q4�w�	��b���
��ȡ���@p�o�{ʉ��w�f�4@�61C�����j��]��5��e?�z��O\9�pq]�Ks@c�Fk[`�����8�/�!^K�z��'E�f��^:m���Cv�<غ�?�=�K�z�`��;1+���h�~Z�M�d?2uk;&.�>��"�HM�
23��s2�U����-e�Aiw5�pVފ����ma,pۨ�����8N��h�����ک|�Ml�4�L>��]�XYE�����X	�I7b��hSĭk���{�=��s0�:Ǉ/#ZyD�s��l�I�#��@M��W�ʂ>.��OcP%�3��Y$�]G�#��mEۧ��������(��g�/�d��ŤC�~[vA��#pi�@��a`����m��Y&�����O)~��s��c^�v�(�E�G�K�;�n՛g!�oF"D!e�;-��cF�D+��?�)ԼG���ƀ�L.Z���ON�#T\�h��y�
���z���ǐzQ�r?��Yn�5a��	p'��)�$�{ɋN�7{�*���!�YvߗA�o��ԎG�%��2^R}� cj�+�T��ݿR*+���y��O:C��=o&C��9t����Ȳ'��ιc���e�,����1��e���f��.ޞM�)���@�X�	GO܉F�.�E7>��9ٰ�:|�HJ��p�?�2������y@�4�u��=�>a&0!�~O���B͈զS�?(�X�&�� ~`�M�:y|�W�1C�Yf���M^E�Ѹ�ezv]���k?\�͏�D�a�q��9_�/>]�ۧ�&BIY�;"	��ѰI�����W6\gK�l��
�b��u�ʏox?G��^vZ;tn�,�I�=��I�kqxľx��D���-x�Abv։�wρŭl��$��o-�b���Z��wl�N���؅T��x���K�X���n-��^�|݇���l|} Mk���xX����ߊZ���Z��~?@�vyFq �*[��S�I�":i�/f��2������FS� �V�  �)G�^<"�v��Ob��V�b�#ȷ6��i
�
��0��Y%�Y?�-�0�r�jP����i���.�������:+�l�7��qH|���ȥ&������1; �|H�Y�b\�I���Opаf�x!�Z�u6�P�[���]h��r���YCo�ne�iS!��:]U\K%�E(IIn�䀉_J%�-�%����B���3;@q�/kU7���^��I���ԟ�����I��'+z���mh�{��x'�,���{�i(�b ޯ�eۏ����V�2Sƚ��.�1��O�Sb(�V����jŏ|��Q����F�qW�c_�
�X�%��c��/o%���E�=d���(��������F���<aO��J#���s�"ڰ��ɞ�-I��@g7ƪ�2B[u�����D��S��}#'�eX|�a/ 
v#��ӱ�4§��(^���濏X��iz�-��3�߳D�� x]��z@Ƴ8H���@ˬ֞
-^}ܖ�(+K��a����q6���c��0|������X�ʾrNJIX���(\1��@XlxVHYEB    3981     4d0��e�o1�j��*�u؅F��f�u���q�#A��_�M�f���hb�'BO-ӧ�$jl�'PG_3C4��{�U��oK��E1JI��Gx4�[9a�:;s�0&�]6�ʛCe΂t.}�-�G�.�v9�O�?��҅�^ոV����*�Y��HO�R�)J܁S
4 �3�&��.��W�Ɯ�1h4��n�!SW�L[����e�9��F�œ��>�7���y�~s��YsTz$t�B��܋!���Ua �r |,7M�-bW��li=[���ox�Ra��s�:r%���6[�����.=�����gm ��\�<V)$���#Jػ+��O���.��y�)n_���K��T�o�H	/���,��ƅ?]��(⢎��������k��LFխP���z���xmo��J�H�F]�6���R �a"�P�?CE�TKv��֪���z�@+m֨�¢�l�k�!1T��.�(��p�����<7��B�䦒���h���j:amH$� ��}�,]�^�8��c�%�/L&������1O:(���hv��z2�ϭ/��j�����&�������:i�0a�i׬�~[�mp���f�;X#��^W�Y��-��v��A���1����N~�O�S����5V��% Z�Q���Ѱ�Q�^bv�Y��o�fn�Ō	"C�qFqb����G�9(�aHw�0�k�l�;�MC�=�ܣ��Q*gﱊh��o��u�(p�
T�\G!�k�	~���2�\�(�)I֐_9ݛ�"�Ț�uƘZB��I-�q�ܜ�E�W�D��\�$@�B�|%�}a��c'<6�<0��d�
�j��0.�V�h=��J�IN��pp�uZ?��?���#�� %P�o�*��F�~�3!��9�^B񘼍O��=ki�����	 ($�)-3r&��i�Ogs�]1>�7^Wڀ]�w@�I�s޵��U�X�H��0���j�+)G� �i F����a7)���[G&���xE~�O��	���Yot\��6AJ����j�[O��7܄&ft��1E�~��3V�]�CB�>�{�}�������
�@1�T���@�h���_m�(WME���̏��ͤ�(��k�EnꘉM������N��V��i�M(�PB����L8�����#X䆁<��c+(Yo����F�!��b}�֌��b�Îцc�!�:�$�x�oh�UAѕs