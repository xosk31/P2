XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���j#O�˄���T������O\:������֯qP����saj!�F�LKUf�]z`6y��!N��N7	�|�X��v���È;:}��=�k��R�$)�-��+hľ�×��5}۲KqHf��i��z�7'��`��`y�Rz��0S��~�޴h{�<O�����a)s<bӥ�Y�f��K��4����W��-8�bGy?=���qN��W��H�8V����a݄q8���b���Mg�ڀ1R�W���
���C��5�?�LX��,Yu0��a��,_$���yjV,������B ��/bVwNE���W�E�SJP��\�1lIIn� Y��O��:d��ԩ/��ݛa��= �Q��Ͳ�6	��i��
Ы�qϸg���=�${��4O�֕��Lts-%{>�.�a�p�����YA�-���ʏ�$���zG1�t��vV�����f-��*Y�������Y��J��sn�1pU�~V��J]����|$����;�||�a J���7�� &�|q�H��C~�Ru�V~mܚ�x�#��0Ų�7�m(`n?�^��4�t�bz!	<~�>���DG���%0=�����K�7�~�̢��? `1W�2A*ӊ�J�/k��Q/ x���oH7}x�m[,ݰ���"&�k ��%1}Z��[в�q��.d��X����Y�RA+PP����X�g1�	�<�j�'�:ȩ��._(�H��$q0T�N�N:�A�V5�w$K��@- C|1����[�6$��_}o��XlxVHYEB    f7fd    20a0=�����9���#v!��� @�j�6������\Py����*H�RY��p��5����4�]��U&*,1��4x��^�M�Y���z�q�rA���!�®w�3���1n�C����SL;�>�b����O��J�~̟^�m��櫙_�g����D,lŻ�r.{�}13TJ@Q0�=�>��H�4
ʺO�8�ˢTc1;���TJ�l�'2�c'�aT��ǐtm*��e��U7f5�t����i��bia��5t"�'U��b/�����ކ�T4�84���Vs��8�@���6�#�sŬ��6.y (�	�3�!=���g�7zm�7]�ԑ���݌ә	���K�jf�j�K�M�^jG���0��L��ܡk��K\m�u����^�U��=�!Z�e߰o2�Ȗ��Ȩx�@�a���I��ƛ�u^��ђ�!��*09���Ŗ.���p�u����t�5���M1uf�/xҟ�z���t)��*u4���޵�����b�V>$+b�eM�f�P�E���T|�[�݈�B|m�9���M�WVf��)�m���⼉��z+���� 
;o���"�^�����VH{�ԛ�����'u{L�3���I'��2J>��wĻ57��;z|4��k���υ�8�����
������6�[�+�]�Hk���|���(q��[�Z��� ��x۲��J�9����wa�Ե��>���z�wh��&�����~2�f��*i�ƲT��?,:A�|-�X\'ցC��� �?�W��K^��CTk=�)�LZ%Tl,��}U�*��Ǩ	0ķ��k���e?
��*�h8��~)g{}{��)��I�¯wՌ���ඁ2� �7�,9�f��.ك̭=ov�C(us�%����R6����� `�t-�Ar�h$��� �WdВ��|���J����3n ���<�%rr�VEij��&e�.�R_����dr$p�O���@��+�c�G�ٛ���\�WT��baH�Dy���RF6�r�����fv�����V�A=M�J&�$�;�㏜��Ku�aUTe��u�)�6�	ݲ���0vș7�cc�{��i���x-`���MNQ�\^����>�6:7�w�{�z؂�z���nt���`��
�1��/�'��{zR�� ��?�զ�+�l�ݝYc7����M�V�$?��}�<�����|k��l���,Q�B�Y>�d�S�-CǥTuS����O��J��h�����
��鉹�<�����+�,pp���T�һG�K�%��g3��E���țx���(�"J���cVҺ�-���a����y��v���:����ϟx����$��q��a?'ǫ"CǺ ��3FX�'��+> �[�`�+W��ੋ��ͫ)��:f6��.�Ca��ݰ]z8�K����Z��B�7~��m�eL�2�������P��_�ӼLɂ��Hl�L��=i�8-��n�¤;���{���?3u��ĩէ�+��ʽ������;�І)� 5b�Ot.��]����q`�ٗ+np>9�Q"���y� �/��E��ڠ�b��}X'�0o���쎙6.�F�医���ꌾL�jj��{ǎ_2f�\�߹�N���+��&U��R9�F<5�Q����+�Q ę><�1|��ø:!'�t��r�@�9���������Ĉ��^~��D�$V04?���N*HϩF�&oȧ	�9p�L�����Kq�ƶ��n�!� �ҏ�������]�N(e?�͔G$iW�h-��&z��E	#C[�z��g���w��O���m4���w҆ڴG�s9J�`���Uqf�w귎�B����ӳ-�\O��)��b2z
��~RT�Xtj��S$ą;��Q%�8���}`K��R�@�χ�~��Du	�{�a���9)���YZ�o:��c�i'8�B|�p�aԋ|��3>�->BX��AUu��i�7����!��s�YJx�"�z]E�z8fa�Э�/��Dy�,�n6w�_�Sb/�`�ͪ��.�>�fڛ�7E������i`ҿ]��HI�� R����++ �&\�k'�@Н���d4W4�����dy�5���0�}��X!������m�g�F,��:�Ø<R��Y�1��[hg/>�l�<\$в��#*�*�B���y���y�����Jڏ2شKI-�ȱG����B:�@�Mw����_���vK>����g�x������_�(��{��0{CYݖ������W��#��Ǐ=Ix��b'i�L�o��G^{�M`)�d�`��gZ����O<-�U��ޣ<TTP��*!y�&�"�c�p��vy Vy-J]�D����\ɁY��3c8��nw��t{�h_�&B�k�A��XdL^_��oJ+s1ƓFA~1�d�ܭ���J���x�hAp%ͪp����c[e�-��J�1$4Y"h�K���ӱ�7w[�>1w���Z� D®����2��>�9�3��oŭ�eJb���.���Gs�zj"VW�[��������\�n�������N Sҟ�4��Z`� .���R�_��N�R`.,(uS��
�Km!~�^�~5�M0���PA��w��|�ݟJl���8ȡV|<%��t~=�CF��/����x���Z�0|nUq�'�#N^�7J�`�rC�4�l�4!�E�õ�b�34��{����Gje���9	�f�C��3���]y	���[�*GHR�K��Ni 3:$2�5%i�JG*��Y"����/�CrA �R�h��Z�NT��L^��&���to�{�㿁,����Ej�F]N x�B��-:�n��\�4�֕�<�b�b)�s��~�t����o����h���$�{�jקd�RO����9���d���&,���E�V-��Ƴ�9Sއ�<�(4~	&2�딃eG�@�r�=�sj���| �Ō��ڑ�!�,���.;�N@���B]����ƭ�xa�><��ޯ����N�F��J�Z����Z��;Ji�!�^
���d�;�.�I[q��m�㛑!G[� ���P���c[�`��,��Xނ�X�^Aƶ'D�+o^�@�N�P�2E�������| \V֍`��<�D�sl(DksBބH�##Ǻ��7�[�W\�ؾ�pAuC��\�|�����`��Ȩ��~�k�;3���d��cQ��~E���ӈ�TZ���}���q�Φ�tAiC��qF���']���nMz�'2	�;o� C��&��ɧ�؉�\F1G6*����}�%�q����_���^��u�z�5n�2�cIRzq����������rL�aK�)>0��V�uR��D�<�A�P���8�$.�7C���|�����IG���rt\;RΆ�̑f��m��|(�qo�d
�cf�PD���ma��j����j�e�B�a3�ZER1��G���/��Շ#�ө��*�kН9aԾ�C�]�p������i��{��k9�u����	������q��(���� �1�zl�%�S����'y>�h� 2��� .�*)�Yi�]���v�%&	����ԝ3����e
��4~K2����8D6덏��=�D��i�L���
�|�}u.�m�#��
�E��/��iz�Π�H9@TF�5"�s/��#�T��|�5]h��B���<�ʪh��ΔQ�-�aN���<f�-1��7!/���l�5��w����f� ���E�S:-c���j��	���4��Bߜ�_?..|�+u(���k)��"�+1�x�>ϗ�C0�΋9w>v-J) * y����2;��>�R�ܵ�F�����di��
��sG@z���c7Dm3ٳ�K�vp��$�7�4Vؼ�.�|1�}R��:��hU��5o%mW$UGF�f�gY�i�1=�����0==�}_W�|���cg�8V�x�� �<A�y�h\L�����MaL���>)J�M��O���ء�1�Q}�X{��� �U\���<"�w��&�Cf}Q+XbE�?�H*�"0���0b�c�I&��O�1�Mnw\	$��x��H���z��h���4S�8߉I�^S��:0#�tC_�qs(pp��ٺ8�}5���P�Ж]�V�>}��ab�_%Z���tկ���o����F�7Z ���sM�ZIL�__�� ~��С�6�Q������eu�J�E�L!Q`��`mR?~�As�ȸ��a��M^�>(P����C�����ޣ��4]Mr�jO�U�h��3X$�"��m����8[Խ����Ks��cS�3�c��aC�A�2�kԔ3�_��kܥJ�~H��G�	"�0��M��%���+c7P��O2-j�VÏ0n+����S@IX��53�v���?��3�]�ؾ*���X�u�S�0��49����0:grw�YC���Bo�$Ϟ���'�48�w�>�X�=ZX?4A�ɜ���gv�tj�Hhw��D84�����N����)�"�K/���5t-�R��:��^���)�I�`���ym�(G�W�����}˨�f6T��"��p�8,�2T;���$�J��^N�Q�6�V����p ��k�{���H�R�$8;s�����~~������eFe�:-Km �&�/�Ԉ�+��9!�������b9��u �8#�+q)7�"t�[��TY���'�X�R޼��sM��T��:��>��En
�^�3�!C /��K1���R����\0���/2�����x��kb����}����c:̉�T^3e� b�o"f[�[a5�<����(�Бo>yV��b�N����J�	膒�t8^1eXB���VHH5D�H&*7����"���F�AE�!s���r,��ǧi�חt��-���$I"��kl���5��(�x���[@�X˭�0����)!��ȯ��r��7��ڙ���e��qF�H*ߎ}lU���Ǎ������fB�к5��A������Z��շ3���2l��ȫ2�bO��S��oMg�5I��Il$��Է.�{8I��n���~DYhS��ΠtM���?�g:��Rp�<�2�4��N�"�JLƏ ˴����ޏ�T؜��z�G�˒Ja϶��=k�D'�$�l"2n*�Iɾ���<����<��-ߴ2����[1���������L �����@�=�M �'�L�Yt��G�k�J>c�cY̱�F9:���7Ez�#��D�R��6��[��x^���/�Ј����oJXP�#ֽ%��c�ܜ'�uYR�����]�ӳ@�W�
'�+���٩�Q��QAa��c�f�Px�V1��S-�E7���(``wE�i�1��k��c��EY�T���u
�����yX�O�����vV�yr���5�T�GVBu�̷E�`d��ha8������(TbM
�����bȞa˷R�#q>�O,��FTkt��e���.�R��1��52W$3��i���E!����OY�<)M��
�vYH^u��ƥm��Im�9Jc�o��c��B,bdBeZ�\���r`�T|��Z"=�:�ߤ>����FL���N�Y���@m$˱Nas!����;?#r{yơ|��3�> tE��8ad�h�\vÉ�dT�%��nP��q�|*�`�(�A���%�����
��Y-����G8����V)w�P]��Fj��_��soU!-����jC&��-�t��{���ۖ��/yF�8s%�od�a�'p? ��A;��T��W� �k]KP���J�<d�OVR��<>�vmYD(�A���K��
B'ܬ�v3��V.�,�47Vҗv*�z��|ė~(cY�bf<u.f��� ��ͰT �ђp<S��m�ףV��GL_�xθ�\�1�.j'�ͷ�f�V9��%�k�U�:��]w���x �h)s*C($�	�C.�ڲ
�]����v��65aH�/�4����_�鲖��K��͚���ӥ��[����Tv��`ͩ�V3F�#�����Xe2� .hx���q��w%씀�_��0~S�\4�^�~��
���%�x�x���|���a�\�OH�$�=��|�|~	���@�Yc�˪��q���������Yz�M������aTMx,�˕��^f3q�g��F���[�)Fp�����,�H2��� ��k�1������B1?�"�
�� 4�Ǯ���/5O�/��
-ڷ��5�ɠO�
�/�n-�%�����3�^%�&�C�·m��y��݃�?�0�V#���fʼ��6c`��p��{����,tWɰ���',<L.���.m;�M��sl�U ��:3�a��fD� ��8�v�-'�$
H^%��t~�<���
5������A8��Q]�mU˃�^׾��6k�xJ��h�v��<���Խ{֫1�����@��`�2 �@�#Y����.�A�4H��R�䍡6�W�y���Iщ=h����N2����C��%M��߈(k,x=���gV���u�E�k�b/�{m����Uf�y�H�.���w�5�9�m�.k�x�����i�)?�����c{�C���P��x0�/����̴2��`#m:��4F{�;�UW� �9^J5��X���82j/�o�|	Xr��0�j&�Z�9����9�M��+�H��Ƚ�;^u���E�||��p��AZ��A6��}��mP�aكA���!#�?6}�Ct5���� �b��^�Vi�[і�b��_e쳩=?.��u��h��ufU�AO��uFt�#.��%��O�2Z��SBmy�4Vg_�&�J��'Ĳ�
��gF��u�!J�j؅%�iV��D��6�#�7l�RI�Y��V��*7��.�ж�w��(R�l�������z2`�����K��P����(����:���,l�o1������k�)ҝh0e���DጪO̘M:W�åsI�<^�\q�2O,�4#���Y�<� �����xf>V��	�v})�X%t��Nqs�7��2�@�����V
��c/ۀ��~��HH��fR���X��k�Tn���t%�Ú��� k��pq?~ �bM�)�|����RU4�	���C 0��^�}�j��g���[E�/�՘�X���~I>x���=$N$V�hm�#u1E!siu��������ȑ4j�� H@����P����c]*���?B��gĿ���G��$�#��sl0{��x��w�[P"���|��BIЩ��mB�鶶��x�Nd�x	4W�ɛ��L�nh ��X5�T��G��k~��>�����CA�V�I��cQT��rǵ4��%tsN	w=t?kM��"Q+q_-a?9h�]Ԥ����LFZ}F���f����^:*ک�zL��lR��?J���]�5�9�Tk��8�A��餪�����,i>^�
����֥%� L�"��
��r�I۝O�\��d/c_oQ�?YߑP�s�HXv1C1�O{�Hmzt�1(���AR+_mN�~T�ʺ�6���������>�]$����[���s��Us@ř�7���g�t���8S�����ں�1:~s�r���>ե�^e�)I�i�pe[��;!12�H9�W8���ܒ㦚����	��,�+<� �Gӣ7۵��;�tm�<W��z�)�l��I�����p�Ժ��)�]�W��d��;��/.�y�DΤZ7��� �8.���f��Q9�W�t���[�C�P��o�gmN�#X<�ڀ<P%�Ru���G�ϩ�攥�~��Ȳ��f�Qb��R�~��\)�=�Q􅶖�����s�~�de����Xz{hA�sj�A~NE$���Z��d�H�X(�q�'�#�cɼͣ�1ri̼A��K�)��Cs_\�S�Ķ�WA}e=�^�S6����Ӌ�ԝ2��o�v������~�[@F<����~|q*�8������	5)u�M��E�����܆���T��Ⱥ����O`D���t��7��P+�*N �ݻ��=���8�����q����q2���h��;(2 �-�	*���Z�~p�
E�W�����c�ؾtͰ��b�9͹���B*C�P���N����X���N+����G�������BQ�i;R����.�>�*ё�<]LB4�Z�I9��Wܒ�u  �]
����Κo���{���DO�d�K�(hG���X���C��C�~�;�����