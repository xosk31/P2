XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��X�!�A�k�a\���7��p<����=�a�LD�#�N��'�[�Ot^B�t�P�q������͜�[��3�`���.*|�]�3�gؽ]��x��o�5��&������,��%f)�#\�hDim�lN)%w߻�T��(��5�Mh`��
d��Y����0�.�(J��9nd����!̗A�_R~�h�fR8ynfQ���0T+����T����`��DV���J����|��O[l�l�-���L�I5ͭ.�Ln�2��
ٗ��&y�PAd�̞��i�OS`�G��Ǉ��U�okhZ�P?��88��-�(����{�E�[4������N�D�9�X��Ħi9�j:9�o�T$f�����C��"I��:����%W��
j�v
@�[�n��R}�O6�b��7B�8)�˓��"����aX=Q��؎��5G���9����:Fc!ܻ�%��6Q{��]������$d���t��qIYv���Q���x�9��mg��[���1S]�i��!��S���k���zk��y�sBMU97T����0��(G����=Z�=R3r��%ܷ�K�dG�4ØA�Ռ�M�T���'�T��Ӯ�EO���pP\f��Q�9]����X��L�	�л�0�v �hs2���?���:,A͑�GƉ�Ah�*���d�dY�,Ո7dW�c���7h�,\�#Y.��k+��u@&|G��c�s�n�Hk����q��W5ֲ$Ñe��D���l��XlxVHYEB    3927     fc0�^�c��{`�F�5� !��x����1�I�Õ���G�9m�Y�`t@��� 4x�������2��^`��uI��i�]����f_�[-ub��~a� >[�1���}=$�k)�a���NW�C�� �H����&%+�����t窧�Cb����g���֮�;��q5��n�>�*������8s�� ~�S-��V���Jas�c-�CLN����04xܲ��#ޛH��Gd$OT!�3V�C!�ut�҃�#a'�h\����	� ��^��ɐԉ�u"cց
���ENC�֒�-(SjN���t�?O�e�||rK&�>�|Ɛ$~w�&MҒ��:�n��^���.���z��=_����Q����F��e�+%�ѺQ�Ӓ)Ie��.s5Ē��$��APNT.�z�D!���7l������kQ��o���,�I5��E^WmD���L��OV�j�0�U���t����J3�l���P�d�9��R�ܬ��O�@�ܗ?x��v���\Ⓙ��qS-�ϰo�w��+䟒�v8S�@M�7�TIC�s'��<�&?�$���;�W�qw���V]�j��9�� �����Fz�'�{�3���f�ʈ�v�m���;�����,��DX�F��f����j�[�"o�Ō1U��p�ݙ�촭�J*��c�{�6�`��؜x�nM��2�d^�_���\��߷�c��r�Tdy��˔��!�*��84��+�7Z��)�M5��hg:z�w�a��m��X1�ҧ��{Eu�Y����S9R��0�ջv�9���
�6�̝�8�o�}Y��h(Jf��fA��Z�H���S�`�����Z]N7�µbG+L.ٓy�0(*=�;7L��o���N{���#Unc`E��1��������Qjr$�rO��IQ"�M��ay|F��:����&��8;
T×y14�"����/y�tSR��V�B�ʡWd\*z�i��r���:�{ 4����V�9�cG�W�;+lp?��>kY@"c��RS����PP&�
���Ta:�Ŗ�Ȋ��f�Q�pİ�"d���A&�#p�,�p�O�A�B�)�x����5	�X?;P'�E���]��.��>�\�w��f�Me�ܑ��e��n�S(i�%�����2�z��v���N��dNC�IL���9Br��>��d��kO>?R#�;��8獝�{ް��Lt,�rJ�7�d0,���V�����@+���7Q%Q��{�`3�ң3G�D�߆���
���H$iQ22s;�1��mr�GH���G<������A똊�b3�+<%�Gk�,G��t%��!gߜ�V٬f��&�����;��<�A=�=\�O+���rA�=;=�>���0���&�-Z��ќ�E�P�7���s�5�������m91t��$wO��w��A7�n2*!o�d.�Y��b��CBp��弮N.��e>0�]�]L'.���âX:��Ůt�d��TQEr�  �7N���Yi�~{j�ӎ[���AN��J�G�)1���;uiH��f����(;�>���8�yO��+��sg?u��.�q�<�*?2��!�&�z�`VO}J9��M����w��W��/oZ��(���k�xq9G�"�󛡖1>����Nqߔ2'��JR��a���Tr6R�(8�`e�?�	�ڮ,)���)ȎQ^������a�w/[�����$݈���$��.�ٸE��ɜi�z�mi̻_� ��t�CP}JľB�;�
\���B+�m�Q5u�,��6봤��/������j�'��P���A�~ڡq�%�6U� ��ڃ �^��,ڗZ��?u�� ��\mK�t$p�y<����$3�_$�c��� p��a@}~�k+�qg1>\]�	ˊ���h�c��@�3�v-�E�~�#
�5�K8����^e��I�9JT����r��*����| c�� %&bx�1�Ka�͸vf��^�t,����Q����~�����f�a��W>���R��݄���]�����fG�u��IΠ�Lݶ�i���]����#=��mO��i��uo~K��ɨ��wC:-+S�*򇪅�f �-A1	t(�	��U,v:+J#5�4���:&�������/�Oz�l�g�5�D�5<%�X8lE9\�P�Q���&6��L	�&�֣Kn�m&^x�������+�ˎ@�m�Q
nOX���?���1��R��٫v;�hT���7�n "�8,_M×�S�A�)[���!ӰqAQ�$~x�xΉ@�^����DǷ��B��Æ=�/��g�:�F�l�RB؋M�T4�o��/eB2�+�{@���K�����i�zcRb�u�(�3U��ȵKu���!���I�y��� ��/ڥȸ�Y8��cB����6��)P���u�'���>F�˰$��4�eQʕE���@\����_rK�}�Hb��z��1eO�>%�j�}�E��5��	�9i"�p������Xדu�fRiʲ#o�b�|�\O�f�J��1����6�#�6c�x��扎Q�ד9��w�Y�T�? �M^�����:��e�����T��?u��
���2Q\�Ü ���,�k���i��O����6)�v#�CG/w��F�c���j�hO�f�6�u늉;`��@��g�ڞ'd���J���A�}Qʣ:�����C&��A��/+ႈ���&ͯ�4�����!V��y0��b��T�Fɗ�E��I�K�H×Ϩ�p�c�9���[��'��A��*{��;V��<C�G�-��{��㚥.�:�[O�'L���Ki���E�%�� K��K�%�VH
z1�%�'³��O4����у��Y��8ᱼ�݈�/���x�j�޵4���U��h�"1?ڗ2�d8�JI�ù��%w�0��}�.�0�7a&)��xБz�����=�0�xW��)�좜H<3��\�ڌ  �Ȇ��#mR��7�m�E���>D//׬dd�'&��<PhY*IA�:�S�Ԭd�/����Y+��!�\k�K.`r��.��Ҥ�GQ�&�� �џ�����%�0	��|66
��KZI����A���N�|�I�7e��:3)C9u���Tq91�~�7v>~'N���Nq�@0��V`�շ��s���a��w6h&c����'��a��O�{���q��c"P�A��SS�t0�c~��?ˡ��s޻� �	B>��X���(����{��M��0'/�Lt��~A��G9H`�S�}ੳ�T�f����dvx�Z��cb�^}�����X�Lh�ps�7 Pwz�*�_U����G�n-q��0�Ō+����Wj4i�f�'0"]�8�_WY�x>d&\�S���w:H���U|-_,�>���e��'ؼ�z  ��0c�#	}FꞴ�8�]<���'z�9ˏ�$��N��(e|e+��@�b#��q)�cMˤQ�����'�/
eD����s1�%���O7˛�z�2X"�'���+�ɋ����?x~�Ko�/��n���~7�_1"KU�?��%�G]���J�ѾGU�a���Yp5U�C����/��C^-ſ��Ł�6x��lk�1_��1 f-�������!��>�n�ź�m(�[`m9��Kf��D讍�6KU7���oǯ���5��Yi�H=N�[g�!n�Lc'��CM�ȝ��L$H,�����mR������q���.���E�d�q�[�'mGgE M�9._��μ.�|#t0;X�����M�&)V�|��^�kٓ��R��+��ޯM�">+F�z����>�y����([|Qm�`D�����[k��7X�n�]a�P:�6�p��2�JԄ;ۊk?���7F]gY* ��߀(�^�g�<������6c{������c?���5�|�i�9
C�n�)w4=�������·�v��Dk �$�(�S��_�"[���{�o9b�