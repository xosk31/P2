XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Af�@�����Ge-#Ғ��v-	kJ8�no�<z����T�B���g��A9Z�Gl�ٮ�0�~'*|h��J���	ה�Y�����u���i��V��(i..e��dxfE�8,A>T@5�Yk�M50/54W���T�.HO�s�S�W��d��'������=N�`3X�V���P>w�q쌩�p�.�G��3l�Tl��ءQ����]&(�+Ū� �E���1�?\�kǄMħ��� u��C�_�������)�j�#��:ʡC�`�H��t(RȌm!�Nש���d�K6�x�����j�m��Њ���VR�}0����=���GW~�&v9�F�~0ȁ� dو���p~��}^V�C�f[���Y.Y@�g��I��qPs�UL�j�G�Yx�PħFa$5�G�J_T3k�z�����N�ANW�N�>�샦�s`T�GI�jt�����@������s�����2����]�4f<�k�M�R7EM���	3V���P{t`��؞�u��z��%Y���Y���zyǟ}�1k��WW�{�N"3�� �����VK�n�@n�W׋�Y�Aq ��oʳ��jSo3��%�iX�Uj����X���#�W�DW�u�%��v h[]��|M��@��-�Y*�f>
\u��]x���%m���^�u��[ڃ[�t�q�iddsZ�z�δk��Fn��wǸ��~	�ь�`M�t��h'ƙM�ȱQ6�;����XlxVHYEB    fa00    2910��Ǘ;B��t��6}��O�C��$h�>@|�95}��@�|	��0'�^����<Ƨ皗�$��cKKN����b+-��%�����v�0~Q�TW�/}�`h������"�C�c3��+��P@l�cTb�m�vw���3`�aw�8�Z\�!��)�.;��;�j�1 S��w6?|�����\��nѬ�u�U�",��=��B�f-ߊ"#�r�� $Ԗ�O
[k��q�
����G�b��p�[6�2��ĻD�{�#٧��^� �hO3�=�v<
�:XԉS&Yk�Τ7߆)�
p8#��;p"�J�o��u9�Q�iM7	�����B����������TNrnY��Gح�;!�m]�Ps�0�|�z�[�|�y����$w�=?��k�תX�y�=D�t�s��M~��6�ub�n?�����8H��\Dͅ�K'���$Wޥ�ނ�ݘ\�>���_�y�0	y��i��H(W�.ׅ����)��P��_�wS��W�ݟ�W��yo^��T���!T�l�.�[Y�Ɨ�E^]_��c��Τl_u7���t��lz������+�I�
$��6X�t�ӏ�z�E�h�����������
���C��4�lX*�����'��e+KjB�I�/3�E�2��1$�ގ;EQN���̫[Yֲ:/��y�{ �y���ۗ?�@�5t��eX��/�n��}��������x�wq�Nm��;��F�v���j�XQk��Q7
��K+�ss�I	T���T+�A���7�1?�4pW���gÚ4($�c{�s��zU��v�q�G�L.%�_(��ě�>�܉��l�r�r����l�;��L�iF�Aޏ'(Ѽ��8%�I�7�C-֠��A� T{�w�L�	n�!(��.0ļ4����[B�$5Ksz����MI�T&���<34�n�eK)�M%&K�)�5�Q�9����F
�%�Y�n��S����E��B���v��0f*�m~��< ܪ4�3�>f]F�_�!� \��Pnk��~�HT� �^�	�3"��Q�늜���{� ��ۡ����FD�C��1L��=�M�TK)[-(��$����)�jFtJ�n��+t��|�j+p-3%'�f��S�B.Ӂ��������m���n|yrc<�uZYG���4l'��!�kb�~���'O,;��]�>N�nwXrP�g5����z5%���(�	��L�?P��ʠ��*�V�m�ݡ�@tk~�������&De�6Ǝ�s��7���ť[t&{TMF�5kzz�7�Z�?=fo�1A�Y�nC�!,��T��>q�I��rc�ާ��#�}�d:L��!�#��ן9����upqKX�8��hi��O;��_�g �܀Ɉ�3�0T�8���xXҳⴿ��ojTb��zL����Gm�V�Bs�CY�0R����Al�Y��1P�4�}�weȀ9��cV����+ߨ(����9()���L(
a���x`z��hn�p&hk�]���'�W��$g(ÊO ��*�Q&��P�R��\@����.�P2+�:�����ת�ʅ��"`��
N�B�%QDUt|
��;�<��ʄ_3�&߱+H�at٠����t���iRV/�;��V?p4|���g���P|��%<�����ֵ��e]�VHey��t��c�vQ��ԋ[z6�^Q��\i��G�\���\�agj���t�&�J�b�����QfU���R��ʸ����&-�]��,~Tx��NW�f/�>�C��������W���#�F%4PX�~d������JC���������7���j?ȭ�1�$�z0��g�\o~4��w������xp�w�d�}��2��0~�;˪���NӸ[t�����i���4����	gP��в3����^��m�hw���M@ѽG��8�p�o���q�o$A��0���R:A����'��dO>�ػS�9˺LWzN;��T5R����Y�8a�VavA��Y8-�᮹}�e۔��g9���#(Z@a^��6�cos	5��0�Zkfd?�֎PJ׼�ᱪ���埯+�i��$m�-�����T�?���5;�W��>Č)���ww̭J��/��h��|��ڨ��3�j��۶����O+�<�GrE���)B�P"���ż���8��q�P�b�o޷9�Ґ���[��|ܧޭܝ����蟪q�u��4_��	8�!^��h�l��u�-���}�"׺u�t�ة���6�� ��$�SN���Ө֖��H�u�*^�֌Ö��j >���@����X��ᢋ@c��hF��9MR�?϶�zyr2A��R�+]kB9RQ�C�iW��a�	�E*��Fp�,`
B���l��H��=D͓�96߻�3�+t���@�j�IB���o�Zַ��i�]�����mE�>�Ո���ӣ�����D�R֏5u�z/eIf/��ћג脬��J���uv@�j�:�}�Ep�����@�҃-.��O���e��]�Ot8�j��h��tX�9:]ur���7A�*��ڦ9�׬Ӂh�DqY�a�L�B=��������7�
�������Nx%��Vǔa�WS�W�I;sS
�@���L���C���b�!�-<c���O�S�.W�u�fZ�z���v�$��I}�n�l]��l
o'i����"�%QAV�'�{�l������t��46h쫸��$/B�º�mn$��_"�o@<��/&C��ϖ���(��i�U8ʞ�'��#��}�u9�=D�''�>��z�>U��ڼ���D�1K+�H����KnQ��}�K9y�w�%DA����ӂ��� Cѕ�L�%��i�ݏFL�h�+�cm�5+�M�,���͇�Ʋϊo�y{��ۢNߊ[���J��"	�{��e��=�������� OC��� }��w$u�lx�p�D*�H�N����q�l��/�ɸr;�'I��m�
�u��W���t�{�@<h?�}2V/o���X��k=����L��V�����UoG��F�w��rA�a]On���1Q�6ÄLE�֚�Ғ�~�o���v�^��G@1dW�B�q�2�(�R�u�,�W��upeZ��hn�P!��2Cr�F{�xjC��3O��@�hNF[����#�J��˚�0J�`�S���}Q�����|�q��k�|��R�ij��t(��T#���T�lؐe�Mx��b��x�jd����{�}f�����fp�� ),j�B����)9�.F�%k'�y�d�� ��u?��7��4}6���`��UcKUy���6��q�&>uS0�-5���h-Ѡtd���+Z��H�B��e/�=�B��|ޤ�3�0�
� 6��-5}�y�2I�p7��B�s��c8�0��׎(}�����4Btm���!SWOG��b�h{h���)�My����`�irpAV*e�N.I�rOߞ�}�ՒJ%�q��8��LS#b �}�lýS�4՘�Y�$��_^-���K�	Y�g�Q0�Ч�+=+��X
p�i���\|�EE/s�����;��w�Ӏ!��|ʝdٙ��&8�M�[�����ߣ�n>`d�K�������d;��(!�������B\܎2B�^2ֱкJq�Gst?V��^=[d����c�Г@ħ>Ǥ��`'#!;�[1B�'�������ډq��i�9��(P��^�(���f��'�)|J�wt�>�:��ˁ,D�:���xA$Rb�����ko��]R�G����%�or��,�u%R�G�3�F�;�O'�������%Vj��$~�dv'68�
v���ߍ��+N׵��I�HO�"LB��d���/�07V���e]�U�/�	#�,N+Ui�
�U/8S�� �$�h�ޗqBG�n�/�ќ�`�\�L���:#.I��k,}�3�8�ZdRO����A0W��jq���1%����]�i�&6��y��' eQƯy����7�)�ˈ	���E���q���ƂMU�ک>�%ǐK1��#Db�-.����q��a(E=p9S��Lɳ:-l�Eܵp/s<S�c���c-���E�0��B�;u�E;��'�ӛdW&�H���S@���R�+�깭yg˅��)K7�2O��h�cQ�4Vc�G<ь��-���|�(4f˝��D���:��S�����sJ�}׿)�aY*�E nK{L�oz\���X�����HѨ���0������H��u��Z4�4�`w�j} o�A��$�i�ͩ��!�[��,�2t�*�Y��39$���p��T_�ʌi̙#Q�x���5nh2���:$���
�I�&�hO�b����k�Q�ǎ�݌�{,N�8�Fn�n���6��IZ	^�}a�k�Y�HW
���d��hUsf0�� ���Y4#����bokh�mh�c�~6�T�8W���7��O���{���p��ĠY0hW�C��-� �i���G���F�,:-π�\d৛�<��v���w�G��?�Ѕ������)�d1�ph ���7�G��3�{���E�b-5��`�,c�{;��f��=]A*,+k����i�_&��Vs3�*�?�ܰ��;��@��gi�`.V�oU�E3G�#4�?/�aN�|�&�yFjH?�*W�}J�|^ywk3�s�e��;-�g�@�\�D�EW�x�E����V�>Bk��k��o�4,sP׆��L� ��	o�u���n�_0�9�#��V�u���YQ6o�����T蔩�sg��Ʃ�����=����ܢ-z�\R���܋����J��gZ�2��i��H;־S�j\�.1Y���ou�� �j�.f�o�B����?}��#�W)/����@8�KE�O\D�v�� �ϳ�T!	~M���4�;A�p�80�EMӜ?G]���z�C��˃����5�ĳ�<���.h�;3"nUa�Yc.mII_��VƧО�Orl�Ҫ1�g*��Kr�>����h����`��ƶ>Ԯ2P簇�vo4�Y �r$jԔ�Q�/��l��s����5X�5���-�'`���{�`�����d P���L|.��:�r����C2��Iys����[�����GE����NX��B�Bp�h7@�~�����KY7�Cz3�ڱ	���%��E[Ĉp�ud37�D�_�7�+���zu,�D�G3_�-F�Z��̍�}���2���,��6^���p�9R�����K���x&�⒳�K������+e��C]��s��!���a�nΙ��
^��0���0����	mgY���G��c�I��ۃ
VI�>+��<�~�%�L��q�l�Za���M��*0�ɂ�o{N�&�L�V�k���7^�����h�j�8m��l��ͫEdjg�:�굅���F�x��0&\-�%	8A�D �]�PTC+eW(�X������o���׋Fy+�[�kM��JN7J�k���hW���Y�&;wꟴQ%�GU��_��0�!^���r�0)���@����ܚ{"p�gb�6��	S�)�$��8�,5�n��t>�` _j	O�]����kؑx�����DM�?sլЧc���`m"B}.���.Z��Y-��ɣk�vN�m`@C�QU�L��Ecl�i �]�����loDm�]֧ڍ�7��-��ܖ�@ܳ�!���Ň-;]Q�=sk����V�ۂ����!63�������WR�<=¨.e;��Q�}�]K�fD�IC���y
q-j
�{Ӓ8)�Y�c����H�UȥY}1iF��o�MB�6�X��E7Sfi��O��ճ8g<Q&y�s�e�?FM�Tn=W[�=Sv�˿�ǜ'k��3C��2irȭ��;�Ƈ:�H5�l��Q�=9q���W�ɇq�A�:�s6����8Ţk��A� ���)9����@qpu/�k� ܋�����*�����#Xn��2~�|�����3��GT�-��1��_�$�����T?���n�y&9�I S2ƶ�y�ߟ	���|�+u��>�	�b�t��b������EV��%���1d3^P���2��	oU��
�zP^�J�.w�^����W`nALĳ�PXg�p�3��%,A�50n'�K�p��K��|`:xy�kB��H��=��waL��'�:�^m�Q1 G����(]�xPt!��������`�:�4��=n?�Z�_�X�W�L=D���e'������Q�I���m���R�-��4>�p75���J�g���q
����S�	�3�<ɯ=�j#_`19�hj��С�]x���8�����3�k:�e�ȳ�������U��P*RK4ec6�\��n2��n�۝~�.�����J��o	��@c���t(Z�{�֬� �!ֿv������b׸��3����?@��/��#��l��<�unC�E��C�w��,%/�ׄԢ>�)�r��u.V/�N���G�]����"��1T���P�b�3�<��&�z_?UJ9�U�qK���>�ȁ)::��3W�=�k���\z�b�o;ОL��:�M?9n�aIn���ܟ{S5�<���+�Di	i�KW �� j���s¹�&�(��zw��?�؏+�����gP����t́N��+�R{](�h�)�,uo[�MD�0}���,)n�0,��{zVy��
f���)���������� ,[$��ڒ����������h�1�W��]!�_�З�Ƽ���	lb��Oq3�@vRK۞�nc�k�-:͍ 7j��G��[>-���3ARv}���o%*lN���:czE F�IdvEF�{�[��L�&���n���31e��(o+rϊM>��%Ĉ���1H�c�[����c[|q�Qw,é�&A�MaSߋ���3&��?�*�����p��]�Rf�^�{��"��V�y0:�"rI4�%���D��sr��h���;kڙ����������Z@�H|ƫ�i�c��� n3�Cq�%�Į���p/v��7�I*�l���>�dϝE�>����	�)�S&<5�Fn<��B��V[������>'@+�1dה��F�+����G~O�!JZ�i�<��y�k0֥#EK�)�!���g���_^[������?|��P�c���$0�҂]�b�'���}�'nG���%i�7�;����jN��.jq��� w�4��d�ߪ��~$����H�G�ǘ�=�g�����I�甫������Q��:_�4�˞����l���i|�&���9��F��P�Kn�w���]�$�UR�lE�q�d�k�;�c�h�^p�FLX�5V>�dJb����0m��3��5+W6+��^8ld 9S9f���̃B����/?!����ʄ(q�WRi�{��\�P�Xس�NvN����w��8IN0p��Ի
�Q��wQS�����5��1r;�_k��q�	�P3�����E�F�z�/�beLwb �".P	��9�����5�Bޒ�:�����ݰ��p�ެ[b��U��x�J�`?�<U����u/�����2�v&#�z�e�ʬ�}��N����u��B�H�ƅ�gΪQ�F3%[��H�;RJCo����p��Ϝηv�r�KS�p��Մ�_ X���T��S��@�ق�ڙ��q�� Ӟ�e!+8;/�4�j��Ӕ1��&G'�������hη��1+$Y:pg}���NN�B%��8�ȹ�����E@��'�ys\�4]j�z��&ő$`�k�m��n��Umh<�?3׍��KW/5�w�j�x6E�s]s���j�.7!�?�h�}h���P�KJi�`���D�J���}��|NE �Fi�sڧ`���e��sD�t����"��Y�Lh!O=H�d�75��學�l��'�!�@J��)!������y����/n<HM�3\rF�9��_]�0�^t*�Ț��ey�ϖ��&j��<�!>�����a�;�}�5��>ƴg��aW]�2S�XcZf%�l�]�{�o��ywb(��|�b���L2�Z�YV�ɨ@���[��h�x�(P／0p��J��������4���YcZ(Z�6W�P ������^fu�����(7�xs7b]�s^��*�!���勨�#��X��G5�� <i������N�N�o�,�ᏖqLC��^�{1�~��	������
�~̝��a�%S���<���ݡ���01�o��x7�m�Mf���)�Ӫj��I������f��~�Z���>���q����RaF�XR�@�z��/���o�!{��.2I~'O��O�tM�z�6�`Y�6r"k���A��#M��v�
]�U�,s	�l��f��5��;q�批/dU�����q�G�F"��z�ī0,��
����6�O��_gCd�XJEw0#��c*��}�?v�R*j��u��ǰ
� �%���p��5J��1c��ER�-��p+�9�xiƞ;�������{��0)��A����>p�R_7]A�^��H�U�
���A����kUKҼ������C,b�m]�,2�W?���1��v*�U\��e,+9�m��;� ���߀�W��x���� P�nȹ���ad�~�Z v '�<c.Q\7�]����p�x6g|2pHbެy9��h�ER�;���
���CǦ��8׼���F�Smb8Zn��W_�*���sZJ ��V$�q���A��?�t���l���Ca�&;���CM�}=�EQ��@
Ғ�g�48 �*j�ꙻ�*����X��c��֑�mm�ږY���q	�_�h�3�]�<b뼙��by�6�*��.)%��Nǁ$���8ȧ�=�5��pIx��$yDk���F):�@,5s/��zIkm���[0�|.]I�������MX-޲oc����3�)p�T*/~U���5�J�Q�Ao���;zG(���:�v߇��? VK�.��N}�H�\߫ �d�c��_iC�l<p���)Ҥ�8�ƕk��\wYeL�Ym�ۍ�bW������0�3��-�N������Q��N�2���O78'24$���:=b�aJ�v�y5�vZ�׫2����-�zӴ��隩]F�aq�Y1A:;�hdxֹ�iCM͕=��ʲg�C4U��bl�?����/�Ɗ����e���iCmG�������	��]�o�IB�y�.� !3o�$~g\/���Q�y��	���M旃+�{�}�
��V܀�{�/�����)�ʡ�!�y�(lwh]�%;�mJ��e5���M��HD�:3w�ӻ��Ӊ?Ю,�s�VlS��7������j��p��U�e,�p�?�ЅB�HQ��s����{]C�?��l	�g2ǡ�i@H
�'኉_�����S5h��v^�*�7%6��������n(M���=�L�X�w����3>B�Ē�+�\���z�hS�c�����ᾸXkVJB�=��#���Ҍ�p���x�k�N��6BX`��l� L�]��Ҿڕ�cM��!������=M�����`�w����{�%`؝�66���[D(6�P���p��f��,�3��@,�@�6v�)>ʁ���
m[���HL�0��E�c��D�����);����'"�Xm)���t�eRlk� ޒ�5��`	f4�-�S�С�Ue�=�N�$�fԽ�#�د�c	/-�{�X�b��+�|��^Z���� ��/q\��^��$2�N\~����A�Ҍ�sz�56SiG�T������&��T�Z�Gwrhձ�s�M���W��ۂ��˿�?n�}�H���Fy�T�=
%3/�'���xT�>��v��R%����0��z�5��ztK�,	���1���/��h��f�[��M��JJ>�~j��cd��ZhŢ�s6ۼ�ns�;��5܈��Zd#j�M�FHʙ^Իd�2�R엾�V�aPv���ѽ���I��}/�{$������dE�!]��\b!��BE�K��S��#0����w��]����cZKNw�OE������L��`�ڥY
j�j�JG��n�7�33��Γ wv,���T8�͗h>,�Kq[\gOa�\C������Nv��R�4��45K� ����!��]�.%.���W��X`N�Y�_���L_��'O��d)5I�,�3�ı-ǤN϶�Ő����Q��٦bá�����V��-{��⾹�"��U:��,V��s�˒���'����U�\������5~�ܿ_��5+�WA�eX's�r%I�MQ�=��^M!`Y�,trt�yp�Sq��vS$��oh��l7v)^������gz�1������2�:R��.��qͨR4>�A�
���2���\:��i9�� ���)#�U���g�GzXlxVHYEB    6184     f80{M��1�8���*�������F)`�~p�5˟��ݪ~x`t��z�~j��cY$+��K����c�)���9zrT�~�# �>�mK6��C��j���2T\����/��[qMJʣ�A��om��9�� O��4zi��lc�f��.56�|r`�V %.yȸ����,`$�t�.�?JD�*e}����^D\��\؉� �O�iC,�
�]�p��c�h(+Eh����G�f�X�5io/�Zd��m�N�#��/�ZH�����O+�`\^esנ��OYA�A�`�$�Y0)��[0��N�,�v2���f8��B����$���bfgR�#t&|�M���Fw�p����uC��3�pʄ��&H%5�h0Aq�Ȩ�����|�F�(�f��C��x{�-f�C�ڙ� @@�d4r-)���#ct�:w�X*��s�*���c]ע�K��'�oc i�핸�C�����4(��6���-��h}�\q1$�kD�hG�i�J��bXA,^����ZIu��5&��%NL�f구瑣o��>��߽Dj:�>�����z �#�P��Y(�+���l
�:ݶ<��=Ҳ��:��a`Z�Er�FO�3���<�7�eB'@��- ��O6��_X�\m�]�3_L}�V���<�R�T�J����Z�3x��N�/�4B�&=緯�R��$��(���ع� �RHR�	�u?e�J �66�1z��-6M�GH�yr-�e��6�5� .�iW�5�~��b��A^n�v����t�<���~�
�x�A-��C�3Y��ε�[3:�� �x=r9<P,�!�/f�-V�.�o$>�1�Y��+c3l�`:��<q���2Yi�G�v�uh���ȟ82�M]1E������c_�;��r-����.�n��kB.F, 0���΅�! �M A�A?���	.������?���7�=�o��wp��8s�azsj�l�yI�`c����ݪڠ��8fuΡ�>��K#A�TGU>&��jۼp+Ӻ���?߁���CNߑZ�F������/߄گ�t�Qg�R�;��Rt�V���kIk;��(pw?.h��gg_tS@0����ĳa��7}y9��
P���M.�31��q��"�T3�����!�Tl�k�%˻a����j�;0}Qc�Y����i��*�<��K正��9�`�3	qR�`M7+��7��+�DV���A�`5k�R�/mx;����h�P��3s`����A��8����F�v"����.D����1�� ��8����B~�- M#�O|`XUg�iH��Al���Ȩ�����A�B��\ s2� LT�p&� �2�u�������[��@ۆͿX���o;E��a�X� �Tc�m�pT�
I��qg�[��I�@8A�>�^�|)C;Y�y^�P������{F�Ih�&Mz&� �d�c�������FYh1���<&M����tx�c_eY�%���W	���E�n y��-��,�w�Q��h^���v�h�����.阿t�������FFk�w_e|R�$!z���d�E��Eޚ�AR�3�uĥ�c��l9Θ����y�0n�� e�~��8�6<�Nϙ3���8\7�]G�n�nM�����ط�z��J�@p%�?�PO1��jq�����X.v"e�l�AF���Ҍ�r�|tS�[5K�r1�M8bBq+!@#�?�9ۯ���Uo�Io�q�����E�t�"�ch�C��*�#u/������dC�3�>���Ƈ"J�������W9��tSH��)����wU�]��!^���[u�V�$mմ*3-?C��v�Rw3&���:�v�,�%S0�oi�Q��CJ7��Ĭ8pK!�YU᧶�"%�`܁��u�*evb� ��2�>�9�~27����{�}q���ӃNg-;�lpff�"�8I��Ն{_��%t߻ı�ra1��뮫����s�S�8��{=�-~L7�%�i��$���qHW�'�L�Υ9�cV��FӬ9?�������0����.a�֝�W�0r�vb�_����=�_˹�op����B>��pV��H�o{l�N+��,��UXS���*bl�`��{���V��U�?��R�#Ӱ}~gw�SǏJRS(VnUDj���6�ca.�+v��T�m�`"21�üwy�^��~���ӏ�!_�%�l�܂�8�gM�OvwU��CmQ�R�%^��Kx��d�D�����l:��B]�J�$X��T�ɦ�7<���>I �^��Si9�F�Ӓ�Yp��҆+�>�t��Ъd-�d|��ja];_�Ǥ���l�ae���I7R�~&D�����8��z������L��7���CY�^,o�P�����ͭ����SF�7��A��^�l��/8�1c5���w��+Ӣ��$}(ؤ�ƞ"��;�3�ʐhPy������e���ğ��9g%�$��4��yR!��o�sf�5����~��ʪH�4<YR����H�
�OK���?í�g�����o��,?w��̱cM���d�yx�pY�b�'qTW�^�Z95 �9$�SI����#�-j��/�k�1U�7q�������q j��MT^ýs@:����b+ftMW^Q��j��9��B3!	�@���l;�m��0�a[g�S[�>�<l8|��5���e�m%�"��V�xח��v�z���.�uL��y�M্q�����U/�P�\ԓm��"���
���_ vI�(�h�u�]�l �F��\��<X�ɦ� ���z�&L;�����{�n6��n��Ӽ�;8�V�R>��I�)R�v��l�ˢT��q�����Hl�3*R
0�` M֛��r�5�]���ZC4
��X=�PX#��V0�iiY�����w�r{���@4\��#�U��nބ�%_��Î#�]>2��Ĝ�/Ԣjm�d+���p�l������V��ײf:���R�%{ �P��~1�t��60�(F���<�����_Y�����λ�ul�O#�H 8�{�#��	�2) G�v���B��,I!9��m�*.�������Pu������3�@af�/@ 2	� �/$-�y=eܔ�im>�ж_�U�G�x$�6o�#��\��j�q��>y�OD��[��=E��ߣ��%��󾌐�hZI!�F�l�9��QfWm!;��%]��E}�����;�����Gl�����h�m�#�P��t�C��p�+9������5�{1Z�!}Rf�xZ�������,�R9}�~�-XB����Հ��
p+Cupb�����Nǳe���I�y}ܐ�x�mI$w�M�卷�f��&;>d�q��N��w�ZS��5�sq����8�/!��P������Xe;M=v���-��ة��[�4�S��0P�u�2p�p�n'����X�xnح���|@�+(�	�S��s4'ڮ��{�B�,B⃩J( �,���CM�;y�)�	�u�	��y����<�k��P��sm�� �d����J%�>5�z�{WU�纝��G�`t��(�^*:�Ǆ�*����јv��Yʟ�P����at�T�|,{�2jlO�@m��<x�Q'�_��+�t ))����1�[Ra��"Wb�9��nj·�m�=�+o�L�m2��F�����"�|k������б/>���u��{ )���%����Q��0��7�&C4[���J�IP�����t�,���+��8[�`9we�Cԝ�bɆ{.QE�N��Y.��)�
�v>[�(Te/���r� �s7�y�^��Ҽu0�3Y��R�K4x���E�9��/,�|4޻��E��7n�#��)���.�J��0�#�E�Aϟ����SdQ�~�/{>
⍛g�9�4l�3�s����h�(���Z��8��g�K�I����� 0�� �@n