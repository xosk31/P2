XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��V��<-�����>�@���C��a�~�{����aEw8�Čծ.�r�f��ۡ���6�e&.��{�?cA��JԶ m���p��ݮ�1���K%�뉳7�m6Y��.����EΞ��&���8�t��?�A�.D��ǹ"Cx����t�U׭TfO�0_&���?�!	E<�d�ٗ�$<=UE� �W�%�3�]D��V�9������������vh����*@|�ژ}����(�ue:v���_�M'�#��t�7�<���t�}x;鰔���}�Z겯���.�5�T��p�A�%����L�A��aAo61�O2|A*���㔤�M,�����	4u[����IƐDx���X��0�aJӷ�G�)47��]z*�3����Q�<v�N�wT�ULz��Z��'�̨�0@�J�ӿ�m���k���?�?�����]|�np�x�T���*HT^�<}//���""U�Z��\vW��gwNƺ���FC젬uy�TʯP;-CE�ܽ1���̄��75��ibB7�k��ְ�������0��χy��Ti�g�߶�:Q�B~_�'ߊ����4�j�O+W�pDD��MZ�U�r��׽(r������ q���L>ւ�k�&�@����s�)�/�`y�A�e]+��2ڨv6$�
��bg5�4ZU����+��T3�<� o����;H��,繃hŎn�E�
�V�%�W��S,�tSDD2�S����d��tE����=�C����
��XlxVHYEB    9732    14d0�36��;��5AI���
�`K����l��VO,�֟׈���~H��q�<��><yI|��mN�qM}x����DD�h��v���BoN�}7��@ 67��P��h�b�	�|��h56���٧C��V!�থ��$v�b6�2a������c���ML��^hta��D�1I2��|5�7��U��G�QN_��sc�� ��μv���d�K�<��ތH7�r[ �>ɐX���Y� Gf^n)�N^�\b� Ez�t�fૠ�}��(WV�̉��{��p����J��KVޑ8YH&)ѱ��ك����|~j"a2d&9�Tg�`\��Me�f�m����F&i��3�у�7�In7|�֑�l�fA�,j�Sv�6���Pɺa�����������#U/�����Z���Y~���O26W�f�Y� <��rGjJ$�^wO���/��1��(��N�ך���W9t�7��
�ˡ��1���#`2��\M����X�\��=��LlJ�"?c��5d�wV���rL�f~��Ћ�њ#ލӶ����0^�G���1o��qF�e��Җd�v��ֵ���i��3J22�i���_�U�](�@4��7�������h�详G�%�{DE��C�ٌ?�5�+$���~��VG"�`�'��_r�8��_T�.���Y�lW, ���VTO���J�a4K�Ӑ,ݟ�n_gy:-���3���CW�V1�pEܢo�L�"#cy橪�m
k�cr �ַ�Bm�]�/_��bxO}��<�����H�&UQ(����ldi*9C�h�%
f~��Z=������Ѧb����E���:��W��;�%}�+��q�Z/ ]-��a�+�o���2D���	�C��k�oU���N�>�����.�3���]{�V��Mv�g1_���}�U�S8	�K�0Z䋀pu ���i���G�=��׻� ��Qq�4��>�)��xv��rV]�=�.fOU5��X����Ƶ���O�>.���c��t�ʐ�S
�^�Ӛ"z����x��� ���߈�M�,�K:0�������+�+tu��Q�
�b_5<P�)�����gLG7p+=U���^��T'�C�f���<fXI�BoƱ���x�@��.H�R K"噺�Ia_���&��Ks ykD,ҠL!*���Յ���+_"J��j�/�<.^d���(6*�L�P/��lO���	f�W�77��3G;��t��\.&d/ ���F���D���A)�C��'����d﹄�uChWY+�-������6)x2}��(�G�9�\�~� �,)��[V��=�D��.����d)�{�n��z��� �$��W�O~��,�H�ʻ	�~��!ѻp�d띤�sE�!ޛ��t�^�%ok�'8�;i��4�z2<���|�^T�����F�j	�1��:݇yY6�j�Q�_J,ͰQf-+w�P&k��<Kn q�)��+�S�\�!��ԟ���w����K�vb���x�0����V�b���m`��7���	����3ק#n�=��Ԋޓ�m0��V��q�9i@J��`���.��HV�{(Y��i�rP���;t�x�?f��8����L�;[p�m��]�q~��,�:y��n�u�� ��d��cy��_s� �UV�D�E�F�u�����c[[�TV���}৛m�c�?r�,�Ҷ�myO	�� ��d�����gL�N{���?]�v	��jr��"8�N�K��^���W�'�;<���|N��b"�	�O
���m !�)��BxG�a�Ta����ߎ=pA�zG�s��:�9�UG9yomq����+�>�?�*� ӇuXj*�v����v\�F&�9����L���!�)�j���%�V�QH��}�Df���z����+}��?)W�VN�2�0�9����&�m�lz�z��D�"uAJdny��(�]*���9���ɓY�M]��W�70�0�>$�7m"\�K��7�VS����5C��"�?��),QiL��ɣa�,���d�I�<����tRm�/=��]]=�^�j�6���	�W��W����41������b��,~R3Hb��cI�	N#\����8j������)��j�d��t�l�&%�	��c��Ax�ߪ����dcp�5T|���Ѩx�b#y�>�tTr�l���1Ƶ��In)��+�4��f�e��C�˙�7L�3,��m�n��K?5��Z&F#K�
��%p�P"��ϴH`�Qk��\���7 t����i$O� ���֗R��R��K�����	48��C+�,��Ͼ���f����iV6�E]�������6Z��$�+��8-�B���\"���|ۃ�Ԉ�e�ꍳ��Bn8�')n.|fo �G��I�Dw���dPC����CW��"���S��ݹ�=�jK%�������6����`�U38���C�7}A�C٦5�����J1l���RřdF�󣏬c�F�O�����ax*��LS*�u`>�kb�4�=
��*���k�����Yw&}�Z��B^߱Nd��tl��&���'{x�2SP5U�_w�*�ֽ��{-��&f2G�ƼOba\t��͵&��E0g��G���<�k�l����0r0C��F߷Ϸ� ן���G������:�ࣶm�1�AB�ͺ���l��Џ���`��+im�?��xt�����jdO~�MԆ��	
ox���j*���X�j�Sx����S;4⥔:t�Y�N̒NOq7ʘ�wq�,b2N˅�����B�����ܿ1�V~a~�L�
�k�.u,�������OV��?1m��ٚ��;C��n�s���S^srxV&���P�ۋx���ҳ�^��G��W����\� ����X�84�����f����I�$��EA�ܘ�a��%t���UW0ͷpE�˖��y����oh��O�2\Iiؐ�|+2R���h��5)�W̿���`
<�Q�R��V��0����|Q���ݖE���&�xI�B=))������Sv�-:ü���R��d��MB��P0dseH"�FwL_�d���^�jĆҷ�?�`g�ƚ �+�����X���b-��6� _��W�|��PߖG{��4e� =���<�r!���N�;f.�������b�ںzQ�H-Y�`Ud�����9����NjΑs��bEy�W"����~�c6�d��E�5�PhZE�o��x�xQ\m�c�h��W]�g��d$a����G^�$o���K:Hv��/V�<�~;��܈\7��Ƒ�"9�p���w>IT�X��I��C�񁳔�Iٰ��%� !Vݘ.I���L&�9�|�y��\��eMV�I���){��ӥ��
�=�o�E"�.�Bz��D��i�nC�͒�0�2m�9��ʔ�0�σJt��{u���SH�*�',O`4��j��~:*�l�(Ī�Y��tϪ����jGx<N�u1�R%z,E�P=���8*�{��堽�|+E�DY��M�Z�䌖��b���i��}���ZUH��������m��њ�')~/�����\�}�iG)�_x�&Ԑ�@[x��R&%z�ioއ�S�@c�yuޏ��_����v�
���^���v�L���<���!]�<�T����k0�k��k�T9I<�C�6:޷���^�'��^��� rM����Z�n���v}�A�q/��)1�t��8���r�{�j��ُ8��O�E �d�p0��	&W:��y#J�K����ݶ">`t�K�L#��h�`Z3u8e!f��U*��²r5Z�aW����
8��2c�؛�b 48�0Í`��	�E�It��I�O��Oo��#���O2�;5���iK7�u���lw�w�=�e�y��K��X��
K"%Y6 .�xR2��,M�
;T�3d�P�1��\�	��yJ
ߵ_�N�k���ރ�͔
�;�`��<$�Б�ө�p�1��DX£��a���:��dP��������#k8�|��r��@��X�kM�ʢ��%�;Q
k�-��eX�R�5)$d���G,��S��m	�A�ܸ#"�I�������{Tt�8��OŴ��5U>�	����LK�7�hi����kk�O�əh[���!g)�>���$�}�P�f��zW���Ƕ�w�5���Z_(莔D���!�I1���f���9�2:X��ܑ��֓$�ga��K	�嬽�����k��ayv��'�胯Đ��ܾ	����}�!�"Sw�!OWO_�uHp$o��u�a�E*�9/���sOTa�_E����r=�Î��+����/q�âW�G��[��7c�k�Y|����U��P$C3{`g����N./���yӸ�4��d��2�\kW��r�b�{�z�bN҈���=��l��N� ����Ķ5\��t4�UVI���~<�g����t�
G��399
��c;�^t�<�m�e���_݋����<k�)vɘ!�[I-'+���SZo��wx=r�_��L�t��A�9�E_k�9�<�ê+����3�X�k�w��?x��P��Q����k�N�w]:GQ�����������������᠋�#���S�m	>y��x���V��T���Y��$\Уe�R�n����3w�ф����&���Tv~[�ހ�Q�m�P��wL`Q�� �����`�Y�6l(��[i������t�@��� ��V��}
������ ���q݊�r[%�`�=��Mʌ/��i؅^�x��pʄ��1� ê/#�ɝY�˜�E@�A����L�B���Oݽ��~��B`�zܢGxa�8��.�H��{��8U0�p�D��%39�����̏���rpJ��������5Y��_��**Ѧ��{\�a���N�!����3����eTa~u����;��J��fT��S�fT2p�� ��K���EN�ө�2�M����/��Hw���QA6�Y�V<��Gw[�"�1p��������,B;�2`���c�_A���w��eui�y��'���	mE����}��h`��a��iGZ��ٗ(�	��{�Kޟ��"��$�x0j0� �גQ��@NUօs�L���M�k�DL��YTb-Q���R�n�u��HO����?CA��!�69y����|��Va�5���GW����1Y����xB���=����kjUz�ﳡ-��DI&�ʭ��Z��nF2��ED?B