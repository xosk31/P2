XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Y���2�1�U�9x��@ntJC�)��I�7��dh3�(	~���N�j�
8��B��pE3����B�㨺�_<�S��,O�B���}��n������;�Ho?���j�O֛Ũ:u���`������Όvpt3�2c�\��KS�5n�0�:��d���}��KJ7C�(�߆Ȍma��[ۦ��C�0�k��O����e%�L��s���.��<�<da^�]ۙ:�!��a��޹����r;�đ*�a�����U1���{��U�KK���(EI��5���	 [A���
h��,��뛓aU�2��0��5������^���b�K�Y�,�r9_�w���;� dE�0��B��B�K?e�s�@��*����>=c��#��I'�K'9�9���4Q�E���p�V���"�<M�a>�B�(K���tT/8j\�J��L#��%��&_�m�f��MĠq��%ws����U�Op��4����,'��'W�/Y��"�3�9 �C�F���T�!��2���Kz��f�Ow���-�mJFܯ�A��3�%+CRHb�I
We,�x��@ɮ����B>������E%p��ĸSW�@��qX-�����x�V�5Ě������J��"<�������lU�x�(�d�eВJ�wb}��ii�B�ӗs��4��W�Y��wNҀ���Pn*�p����V���ᬧ��E��"G��YM���yg1
 9��@΅��re�`e��� �(����&�XlxVHYEB    160d     7d0�X���ƾ�*�0���c\��-�2�Z�^��%$��2�D�;$o2�g�6�сRܔE�7<�t?����F͖��bY��-�`���KV��.��D�$w��1��w,\��7<��Ci�v�
ڶoj	��2;3:��rY�ل �L�t-�jd�&�Us�i�Q�Aʮ�.�E�p�4q/,zܚ�P��5\��_F�y�w�60�a�����0�1�-�� ��/:�kɘ��>�QېH��8}���a?�$�6������1Aw`��[
yQ�RG3e�?������/�֋CH}�ls*)8![J=G?Dq5�C���)U��r���F!����O�eыW�r����S��I��`��`Z%#��̙?Η�����Ԅ�vXSaL��?-�!%"�L�;pCũ�A:�L]ڀ��~m����K�Y��.az���^��t:F���ա g�k#�n�C���Z��B�Jb��H�����,D�Kp�2sg�1;��͞-��s�b�4pX�z�6���I�=��Mz}�x�ךW��p���(�g<��d@�[+�0���&U�+_��mͭ� �ј��c�Q튧�B�#}W�?|Q%��:S�O�B�/yJۨѝ;��wɭ��Y�d�����beo=��@f5OrV�1�d)�_� Iɾ?��T�s��T5�8�Q(R2: f0�˻����S�D��x�3XsUFA�i����1����ʑ$J�R?ÂhMVa�K�$R������k4�����*g��]_�ۤ�!Hu)�k��-��x7C7���.2S���@<a����H�K0`��ʌ��:Gh����K-4���?�M!��-�`�+�Bl�)J�ʣ@��m�XW��T�9	��Dw� ˙�a�Y�[h�Q������v?��X^t������(�YW�Ø�8���uv�B zaIiޅ0�'�[�ig��L�e�`>-%�f�+�k�J���vo��&��������vV�ũ_8T;��9#z��\h���X8`[y�:�|�>��w6^c���S}z��P��*[l�V��w�A�?��!1�ey �pמ���w�A�ld%���u���Q��̿�<���$��<}O�I�뚍�����,�I������U���(���7Y\��Ԕ}��!v���XX�ۓ%�곔]?���y'z�"-���=�9��,,����+�m{_d���� p���sr�dU��2��m��B�ڿ��M�Oc2!��V�HE,�O�ǒ���_4��4͙����y�¹����ERk��9n�?��3�8ZlF�nLa��{��4Z�5�.��^N<�F�����V-H�HVZ�(�!|�p�b�ǭ�eq�?�����Wޣ6�@΂u#���%rq�ep��x��A��}SZ��߽�o����7��CHﺚ�À/��xF��'Iȹ�2�
+"}#V�)8�����ʖ�*x���P�Y����������1_1�>;���Nq�o`U��y+��o$��+"2��рl?:�rgX%w�>>��h���'�wv���0�d�@��r�J��6-�}���8�[��q�5�'r ��T�~����=�0�@x��T��U�%�o�oG�'�+���n�I�Wo�bѭ�י+�|�:�Է\��^%n�m:n�66b���K��R�cp���V�V�uC���j&jcI#�6\ٟ<�J��Gޟ������=�nlO-tgO-?/!�}[w�߼ݓ�*�]@9ɹ���(���#��.�#����Ρw����4lXo �=����mn���w�!8u�.��g�G5��K�^�&S: �}�B��	k=r��!�4��քaw����x�Zz���N!�
�������a��{��䚥��3�����§hl�#�K����͝��Y��4�fh�U��� �&���ؾli���7d�4� �_;x���K��Y��~