XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��d�@j�((?򜡷�):��@�(ٕt�9V���i�a��_�X�la��KUL`�d1���Q�-H��>�J������_l�v&��1��ׁ�����g�  .��ݨa���Z�$H�����"�	;�uY�m���4h�aj��UZ� n#Z|$��=o�
E0�����������ܠ0���_WR�^�"�����bxg����%����򥷵2G�<��n�����~b�d+��0Vd����߬�=�:c��`��<ILSvw���۵a�����j�y�1� 1پ:�^��ّ���g ��S�*��k%�{��FXE��i���.��5!eiP��E_�t�/sj�6��cϞ�|�O���΀Ǖb��z�b�t*N�L�Q��T�����4��#�=�$�������%�G��y��R�c�np�hpeC����9�%��Tc�鏫�T #f�W,����@cd�԰d�9�������ދ����\v������]�=U���X��RB�Nb��������҃��b��������)��`�5�M�h�?y�a���̽��ۥv��c��Q<i��9>�ʜ�)z��b��5��ϖ���i_f����l��:�B�'en�"{����s7QC����A�'�N��p/�����w����.��1�v�����ѽ����)�AD>w�����0T�2�	xHEgC���A�ы^�� K�9T	�Z�_�9iXlxVHYEB    1a5b     890�@>����;LS0,K�~:Y�>�n�\�Ю�U����ˣ�Hm���/)�?�l��V��3D��!�<�ܪX���83�kLNݗ������O��r=%��I9!���o,�Ŏ�F'^������е&��Py�F�" �!lt�W�^�ǔ����LtEzl�ܚ���F�?�ڃ8X􉧗<k�0l�:>{�F �?���q��0�'M��c�+�ׇ��5E1�s�ou�cv����μ�޿�ű4wa�ƕ�m�����-��Tg^���Y��Gz��z�13���x�N�����Bt�$���ynz�N����n�B�l��$��?,M.�&)q�����,�*�5��_'g�~����N%Fl���wb��w���Mڄ��[��ġ�8oa|Y|�+<���� ��xZ՗��8r~���#�nn3��b�|06�0�����7����*т�+�����9�ؑ�,�)�|>�a�	��a��b�i���9�br�>��^)�|��
��Kq�m����t�����p�#Aa�Y�x���n�6�n��y��Y�E�m��4��E[��b��%�-*.�
������^�s�EZ5צ/�d*D/B(HQ X��䇿�񳚴`+c8�cV���^?ŀ�ϪI���Eh��Eͷ��3ۘ����q�����i��⬤�;ϢC���֘�ܗ"�%�ƍ�"�d^;�VKz74�C�Lb�
Ŷ9ÀG��C!�i��,&�k�=e�[�ԟ��f�"-��ߒߘ��\�!�]�d�$��:���x�B����7:�M������ 1/;-I�b�j	r�ڑ�yYR�b�uJޭ'�!��h|��`bf��7���c���˝o<�[�����[e��xKL�DVA@:�N%$Jg0�b�Ǒ��-G�Ĵ^��09����`V:�"%R<����Τ�|*���}��8� �������N����������LYE^�\@�Nx?��ez�{I��4�x�zS�Y����
���AݎAޠI�J�w����_�W
"���T��7V�ŚX�t�դ�C*u�����x����}w�rUo�B"G����w#�AH}+C�I5*��t�����L�*���]�`�8O�g�nEۯ|�$���9��j
H⧂���d!��fuS��G
�	���> �y[��q���K�!�s��A�ʟȞ|WSr`����̶�A����H���ڌ#���&�o?�>60�Ω�z;9�I�\�lT۬y�	����g��ё��r�r-����d����l�<���� ��`9׭i�t`댢�&����a����*�H�
	�,6��;˶��+�����ov����?�K�%���ƼN�O0�k
 Vd���ߓ�.�����c1��t��K�rG;д�3qq>/sM���>|�_�I��s���S����2���>t/�J #XN��ߪ��q�;�K�r����<���*�ak|���|�j]�泱�zl��GU�iU��L��� tȓ�����:1|�l�v�w��	��l��ń�6�5i>��6�~#*���l+�Pi�`D��|�f��u�Uɴ��+�K�#��"��'��!�|���N�7��Tg0h�]�L�;o�������M�1^���L����%w%d{�6�fY�Ԋ�@����x�lX�،��G�-zdw�+g�kFEPY�@3��A��T_=�t{'����{u�\v��2�����JN���8�a�|�'�<���#0`�aD�,f#�5���R�9*\dz�`_|4�����Yib�qW�;`�I�&�[	^}V���QKӃO�,�ҋ�Y�,D㧿ź��֌��X;�������.%iu@/u�1�����/+(���Ϗ�0�Q�欉 �r���cd��2�/��b��g�MG1������| �\�O�Q���j#&����6`駗6π'�\��H.�g���Qh�a���$"��1\����k��]�[�f�C�SCBsm�M��Z�c�1$�[�m�j��P�A��O�����-j�����*65��&x:� E���y�Z�̰;�S� � �`4�E�˔{�p[q�
֓d�:� �9��J�>��g
�-���Xa�Cħʸ�yw�nX:}�J���
5�BZ���{���t�oYU�|-Iy�]y��