XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��U�;�2��د8'��[��ïO��3�� Ũ����F�(c�oA>'WҬ���&��	��R�gW�9\����6'�Q�X��K��d�
��ũ���:T�Cߡ<P)�:��ry�vm.�K��	�iHaHY��Z�t�T���++�B]FM���9)Dd��l�*�8�� C���g��&���MV��w�@��U0�Ӽ�@�D�P��	�L���6SJ_������L�1j��@5��$0=��զ[L*��窝3k[m��$�Eۓ���/}p�}^1�����=��K)+9�G}�?�pv�A�
�N-nO�en��{�LF�[���
`�̌�p��np�HR�1���]+���b��et}�6��ꢨk��8N��U1��T�kπ�{�u�'����������x�é�"X� ��jV��̟fm0��6#����T�l��9S6 �-2V+�=��H�r�:������8�~��h+����~1��荃(��M��cR����ů��.�8H�i�����J��q�+5�|��}/��Q��׿��� ��A��^h'��������>��0��e�,�<w8��t��j�6��q�����V�[&�q�e-˘vY B+��~W���+�=�>�B?�2���⎇}+"�-pa�R��`�4t��:��Ͼ���R�q�5�M��ULK;;��l�&�p�9Dg���M<K��DX���.�:$5���Z}�?A�P�(����j��q�(!>C��	 ނ��1sX �l�j�XlxVHYEB    b631    1a00>����� �H�>sE�U����v��}�������=��з�s� �Pos�ꂶ�F=D��& ��,y��`K�a ]��Q�T�df��d�l��4��݌]yl*�Y������g,[$�����a���c/�R�D%{�QL���e���Zy��3#�w󴨢IIJ�J6�8R;{�I\�_"�"���z��(u���27���Vc7G�H�H��N|s�)�zh,L�`Ũd;"pFt�t�=���ltR���]�rRŏ�#�# �>�+}�5���)�9��q�RVu��*87�e���ΝȂ�ѯZ��.E���5L+�CME�c�v��V�H�W�߾�ן����9+
�?�g�%Lo�{�q���f �`?��R�y������k/�pR]Όy�,�`�!>I|�Q�w�����;���G��PkՙGz��h&a֗�i(5g`����~~'
	�[���� >j�diN��cr�� $��������;�ap�y�j��v�q�'�r֑
�Q�/`�?�e��b�[�aֱ���Q�������`���tr�H|�6��q7�}v�G �+�������¿H?�x�#tK6�(I[�a�'���B��qڙ�����Т$�P r8T�ߺ�5�G�Ï���a�HGv*]ޗ������Q|��1X�Z��Q�Π�vV��f5�B�(�$(^�4O�K���Q���܄�I�b�6W0vJ��iK!U]B-�J'� �;Y����|�o%%��̔l k���O�}��e�ͱE_�H��1�Q�h�6���K�+;�}� Tj_��� 2��(@���T�r�!��މ*�?\KR������m/�쳵?��.Nh�u�����_^
 �>�N���K��<�x��������H�����������}C����:��W�u$8o�q���v��'y
�n���`y��O�Ԋ�:Dv�XFuU�������~r���8�I#�V��#�OD��%�<�5�����)ԳD]'%n0���D����s䠤��z�f�~FF!�E�m>ى��۲�G��P�K���^w9i��e���x�C(���þ��B
���6�"��3���\��,��	.@��ګ[�¹3��Ǐ(�IǤ~B��C�D�ǌ�ѓ7��(���Ai@þ�H��s��ٲ���>��T�«�6��|�C}�x�H�r'�j*Q^��x���9��r�����3���G��D`���È�Ra}v~�N�f�l�7j��r�6_�\5Z����Z1\��MH�~|;���Dt��S�\�7e�L<��R�n�(:,�>���Q��rrBp�7!ܭ4�߀�p��O­�܍R6��{�ǥۀ��<�H�&U*�.�V!�P�FT���[��@v������h~�sú@\�#r��������(�+��`������U���>�mNEo菟�|�`rӟ����{�+��.�ެ��'��spt²7��^;�:K��Gv�6x׌�/���b�&�$��g�};��F�Y���l�q���E#����H�i߿@ꂴon�[`	eԂ��I��LH{�g����|�D���#*N8�Z�Y��b}؋��-������	����)@����{T�QOr��{UD$� ����$[<Sgu�^ӂ�J����6sΌu�(�+wꑎ��ۦS�f9�HJ����>�նg���ce�=$���o��,���<�9�2/0����G N�k�|�:�>�j��Դ����5��xf��{ѣ�Q��G�%b�_l:��Y�b#�;��F�Z�V'1��A��z88�lwP�w�L�/@�9�i$��qBy�Pz�����,��7�8�V
54c8��pY�W���k�9��s�U��	r�S+,ĺm�_��{�8�ޤ�$�>Ƃ%��z�H^��`�����`�1���!�@��;Y��\6(.SCa���2�Ϲh�Z�)�~����PI؂�\dp�sb� oE��y=;�����'��8l^}\t�ica��-%r������~�ɠ�.�#��`グ������Vf��q�W�{���9�#�+	r@RoUX�蒍籂�BP�҅
Tn2���y �<������w�N&�s��g@tsd߯`�x��Ҕ-CD��M� �$�{���&��a��[�6V:`ڲ\��3zo�(pU��h�b=z����q�ן9ܙ�rN���1�ű�� �9>�.Q�s ���}�Ix��
��m��elO�?�x�� �x<���L.�YSϼ?�,��5�{�ߙ��1�&h��g��jr��ξO,D�|K�g�X��p�z�Њ��k�њe�ni�I��k�u��E��h?��"�w[���T5��&�3.�x"Γ��^�|�%�,�-�K���VmV�"R�<��?���e������Mb��Xmtͧ��߱ޥ}P���s1�>����2�5_3V�I�c24��E�Z�~F}OY^��ӘN�W�gZ����"�U�H%A�ˢꩮ�[S�y�c�ݸ��q���SZJ���`>=G �r+��f~h�*k�!��M徳���B#
i�ǈ����!Y�������WTS��`��ԩ�w@Vn��d����`	�Zg��˵����u�5�S|�0h�_�5���x�P�A�.���ՠ�̻q�6�bǜ�'&��G��!�ȃ,Z,���
&�0��=/�K�\��@��BqT*/��iD�{�����L�tOFK�*u=�V�x���	����7ɅW>Ɠ���p�=yJ�e�=~��(�D���[[y�_c�%��B-��n�c����J�+(A �x[+\�脝�������]�P&�z�=#���Gu�)��ãH�(��OƏd�g��s��ȸ�"OKRz�S4�o��.ػ�.Z�/�_�*��IX�Y滟J=���b���$}A��@�U>���dv�Jʣ"]��������s
�sK��|�沄�ބq�Aݣ�����3e�ǋ�G.p�,D���z���P�N�h�L���-p�j�̲_��0ވ}������ڝ��B�s��V>3�3�
~�����(?P�!C�V���L�����b\O�?4�Zn�����(���q��;t'uֳj�Ed�K�v���^�!W��M?(�tw֍W��k������5g�y�7]�+j��nΏ��X�.�QA����ӏZѻ�vlS�>� �;ָ�m�[?�]�T$�u�H�mk�Ҷ�lm�o���g��wV2���Y�S�;5��몎�e�*H SoL��.��V_1n�t*(���d��
oFA.��'�yJ8>�s�F�)ku�Ħ� r���8	�C)F�J��ؿ�����m��Р@��Y��ۛ�5$�U�A�\��ޥ~������Cx@���ğ�mg����~�K
�K�>���NY��o�=�`^B�ԛ�N��E{i�(ڃcK@�fo��3�/S����WR�(�RO���?�$.nhb;{D����)��ˢS��/௅��F�#���ބ�c#˳��|�����?��j�-�@	�EXВo����[�)���ՙO��jB����@��8�n꽂k?��$4p��P��'$��7gk\�z��/[lz/�k�*�
Y]w��C;����"-�c.�9�'� �e�-𣬝֑�!S�Z�g�����I���Wr#n������7W��)�c������B��*<�+�z����U�LXg^q>R���"l��Q[V�Q��Nӧ��S���
;�����:J�bqxa�a	�o<�a���Gp�FL�c�d�iB�b�ֻ� M����ɩ�l��j��� *qB9��qy4F%w�;
�zp�J��%��4�}�"E=�d�B��Mx��&ƾZL��B�w}�K��ЈԴ�E�;�N���L��V2��ْӧ@g�$�*Q�Cp롹d�3�����&�1v�&:߃1^f��o[H;`.L�$!x)F�{�<�9�~
|�O�w��vxl=#~�"�0����lҸ1�0����L��̉#�ϸ��nyX1�~�1a�"b]I16�縷���3�o��?�=⡄���QS�:�:4�����j��G�ř�z�Z~~6��fxY4y��P��;����j������ #�=�l�����G���5�C]��$�{��d�(��� �2Lo��d��d�AHy�e���Eop���!1�\���E/�gp%S^�?U�(D�H�^��0i�����v_�PGT( �T
����L���_4�Ӑ�7�8���������;�W����ޤ�x�?�l�d����Y���|������x����EN�(�e&I�I+jQ'�j��G�3O!Դ}E�%܊C	Rð����C���<��6����z�6Z�=��Wo�/��e8ۓ ������r�".\���G�,�v~��ڋ�����eF�����zs�fK;�8�<g�|�	EPW�F���BDG�ӎ΄�i1P������P\��Jz?_�;���p<��� �a��&].����ܨ?l;�-�8	�Vc�Z}�̃��:�}QO�!i�X��4j�~��
-(������jl�}ē��v�űx��>໲�fN(Y�*%gJE���F��4E>R%����e��px����xU�ֳ�&|�[��5Fc�����LΟ, �W�5<d�eBr^�k+��.��/<�0�g����X�\a@�6!Ě����vP5A��xmz��㠢�������"���ah�E��8Ux���a�?��>CƆ�q[Dͯǿ�䂣\'��lE>\�%~�t)�lJ i9�xӦx�m+'0m�;���> ��s����J�q G	��YHo�R�VpE�3&�yǮ�Q׀�"n<mO��'u�^�o{��u��ޛװA��Z. ��X��oɼ �Z/�o�(9��,:IRPK@��o��8K<u������e5��(����n�ʩ�R�xnQh�r�Ǐ5�&:�������S���C�?���XA�Qu�2�+�8B����>�D��-�&a/��c��Q���(ϻXyr>'B�%j"Jtx0�{�h��թL�l����F�3�?�L�����n�y}��H�i<���t[V�:����G�ӏб"������z���WފI�6T*�:Z����j�F-'%>ϩ5�������t	�_�9i��K��p�8�Bm���i�`���`7nOx�C��h�E}ȃ]�oɷ<[�/'�q��?��)�6�(���t-i�V�m�]��|��hX
|��Cj뱕�����+�a�,�Ky��mj��@�hʧ�=S�"��	8�V��̓�I�D �й1ܲ�C�,����J����Z���(�κ��瞵���3�E��R럳�+�`������ k�4곾�,�JoT����jP��DW����=�6s#r_e�_F����1��]��{�J�Z�	���~�����n������n��[qb8��n���J�k�[ eY	ۍ*
��q�Z������@��A[)���̔� �ה��V_��K��8�c�6h#4��iT2�-�4��J�طj�s�������rQ�K�����)6�����G@a۔B�)1��@P��9^�WDƁ
���
��O�Q�z�`�x�@Fd�n ��Naϓ��j�9 �.�j��A��&���V�x�	ma!��ϰ��y+M�ɐ���@�ހ{�ꮆ�p�m��,z�����m�oxZ��uI��S�Tt�Z��T�V.S�{�Dy�y$�up��y�,�&��d&�z����?��0�r�c�!O�����3�b����8C(x t]B?hϔ6SX�l�� yc��]��s���_�������c>�g�fD�3�rQH+���j�U���@3�0��������E��h���<�
2J|�t�4t@�w~�ڑ�ی2ܣ��oQje�
���RYF�9� �	� ��A\N��*4�1O���׆U��Ty�I=Q�����Ri���L�[v�����N�k�q��T�Bγ�R~�+n�\�A����Ah�����P��Yh �yH���O�p]|��0 {oQ˘��A޶3�NI��l��|�_F��d�<�ZS�'�+�ա�-*R���z��v��q?#n�?�  �2��{�0��N������Qv*��5'w���^F �Q�__W����2�@'��r+�����d�4���<���k��Nb��i#�+�'Dd���Rt:Կ�?д�Z&�˚e�ʳQv1;(�$&���B���������"�?�UJ9���E�s���	����_�X���k�/}z��K���Y�6%"<̈��E�h�>��.���!:��<4�6����ՠ2w˂,�(����/N��t�W�"�d95Ig��a�1G0{Ɗ ۡ�#����	ʶ`nhƞ�֔/��muAL[����=뿘�=}��Վ��?���� [���5f5|rSr�+�8����	!W��"K�_du���� �
��
y)�/,��ژ�;�σ��t�S��h�X?T�	�Ow?zz�	�tG�����>�ʫF�߬,�\$>WAX}�ƒ���X���m| =^C�L�.�ǆ�����bM8ջ?��|Drx��