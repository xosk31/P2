XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Bw�ݛ48Iy܋�?�+�ٽQ��4hj{/;*A��������-QB%��v⸵ա�����,�vB�`s؀��ǋ.z��m��aE�RaZc��﫛���)w_�Hd�i*V_�w�H�
4���W)�!��4q-!?���Fe���L6/�D�'��4=_�]��a�`4y�UF��pH=�s���q�"����߫b/�'0C��5��m���{:��v��e~��za8M�-^"�u�y�$��.c?�%l�~�,w,x�M�H���B������j%��(S��W^3�����Y��M��1��<��[�U�Z�a�y՜��jW�p�e(��n0j�!��l���a֗)��h��)v�8u,��O���z˶h�r��SFw����%�"�h�5�~\$�����������jSCP�!k^*����q�Mz��5~�tS�R=
��m�핈�ZW�th90ݮ����TD�
�]�-�(��}���9:������c�>ݣc��xw�h_��ҍ9*H`��;�>F��	������Ĵ[R����J�~��&T�F-S<	��|�b�͋S��DО����E��=�%�"����ȕ����k��_>{1����T�Y����@edG�a#p�J\�����5(�]�:~�˞F�E.���������ؚ�S�����(�t�8��<���#�e�2�_�U��y荿%����,X�?U���#lYW!�0c���ð&�x&ЍRS�5�e̸3�#�#��XlxVHYEB    5694    1290�
���N�Q�<���}�_|H%'<��5kª�J:��p�@������t�.�7\�eFr��5e���vz�jZ�GLT�R�S�,@&!����@Z��6�3�P�4�!���L5�E_���c�;�ԉ����]��D!|7�%�������̉f5w���?���Ɛ��u�W�S�d�!�]�?�N5eg�_�}��⻡Nc �����V��ǲ����S@�TI���a�G�E�?���l�S΅��Huq��+�2O�ϔ'�k�F��[DM�:�d'�T�Q�<^.װ���}��=��{oׅ��z�z�������8��� r� �����7��c?O�Φ�����S	�DC7��"�T��u,w�	�K�kЁh���� o�i;����/4瑟^�����hރ�C�^ �R�j����p���Z�7{�i��IT�g�)aW
�v������Q2˩{�&�
W����[�08"U�`��T e�@ҿ�N�Że?B�@N����D�j�gY/�-W��]�}�]�[�4��<��F���d���[B�B�ӧ�1 �CqẲc�`,r�O���e���Y�ԙ�Ew�%-�����	/�1�جͭ��
xP�4L�`�	.g���M
,�%�B�Q~������a����ߟ��0�ͻ�{1w^������|����q/b���.p��&���s=ӈ%��s'�M���a���_�\�uX��%�ı{�v��W�lG�3��ˍ�{�J��b�y�cbp��/q	X5��=}�_p5h�,M̞�B<��m����pQ'�G��wఠb�w��>PV�N
'�F)!!ӷs�[���}�1��Qz�4)�f�!��iW��,*Z)IG���6����U=g��V7�������,{<�!��<Q?+|%<�c�
]��&^��K8{hu匜n� _���Yg�S��%�W�;��I35�3��U���zS�<_R)���')d�b������M��~��JA(Κ��dؽ ��Y��TNW6aSrJ���ŭ��u/#���6Z����	Ý�x�`n�PEġiC�ˆQ�Y���u�d$u����,1�-��W�NL��U�>���di����~灃����i (
!�����#
�0MW\�\���![�PA�9|��8�솬\�e2�|e�C\�l-CW�'7C��{5)��=�Ix��k_�rj��'�Y����ˤ`=I����A�l'͹���2����\;*f"{����=j�qT���9܏C;����}��$U������;�e��y�U	ͣ�T����4��~��`��
_X�K�'���	��YLht>�����~��WKX"�Q%=�ZF
�<�qM���p��XNrF��6�k�{cX����(T��3�x�:R/:�<\�7�j���jh�B�g���K]���)�y"���}e�瘒h�Y%x������w���(�Z ���	��K$>àa�9�f�Я��-����y{�^>"��t2�j�n/���aBti
���~��U\юm?S!v�$5���N>���cx̴P�~��}���G�A}�ut�Xϋ�}�n���D��p�D?9t��CI�K�Es/l҉;
U.;a����:LC��f��L"C˄,dAD���#g!�CI��hn�����%��!ZR�5+�_^%�*�փ��C�`��t�?
�w��D�H#UD�\k#��Mj�K��X6��	�5����/�����^�.a��Gf�R���p�M�t	�3�����DP���x�o��O�[�����Uƪ� E�B|`MO3�Y���a�oI��8X�md�7���m�yn͈ݥ���GVM�a��B�M���Q��!A����5�V���Vl������*i�����(f�p~��T�_V��1ϻ5��Ԇ-�僆"qq����W�R�^ ��'[qC�r�&~	��}�G\��6KLa�����{���_��T=�Y�e�1��0��Yӽ��b��z���C���i0����p�E����׺/�h��y�ضzU�\N�A`�������+��`���x��[� '���mi���g�K�6�����R���J>����A^�[E��]�J^��Ef�!�<�A�-�����Si��/�W�<����t�{4�;����2VH���+#�0�p��k��[��=@B>�͔y�,�Q�]8���-�O�;��~�2p�2q7t�NiF���<��ޫO�-X�������::P����T0�~r�!���Jx���h��lSRCϱP,��dXd��W�,�*'y���D�my��-�Y��/�
K2��O��"��3|�3 oL0[Df�5o���Pw���f򒟁��E���7��J��,���7]7����/���߈���H޽4�1�i��߯	��f(�g���6�A֋�ݺ���%>��}�yD�Q�3�09�D9��D��⨵xi9�o{�I��,�Ǆ]����aL?t�'e�0��s�m<�.����6��]���;��L��}��/��TS���=�����&�|�	�{D���fy��s.�	J��I؊��X�>�#w�V0�<���W�X���-YD�":u]R�4���8Āx���� ��Y�s�Ḓ�,���bάy���3�-���{j�B|nI:�b������"Pǅ9r��D�L��z#���5@G+�yͨ�H4X�9H�T��<�]}���#1Q[�M��`��3���pA� ���97ڥ-���/�n���7��$՗��j�[;�\��2�P(�U��s�Ip#gp=�F�އ�`��ʖ���f��3�\�W5+I��3�J�7t.���^rg=m�U~x2q���xn��P��R�\�'��x��j�v��F�s	W+�ER�Be ?���PC�GpQB��\��b���׌6!�wx���Tj%�	��Y�Uej�-�2�瘝>e#���]��vk�Z�`$$SJS+U�� <��v~�F���^��;ɳ���S`]cj�S>A�W�1�8��h�W�F�k��EC
��{��6O��["���-�g�&�D0�`�"��12XѨ�$� >�����<�L�Eo
,�"O�[IqpG����:�`L9�����{^ݮ|��.��{�)�d�Hz�%�d �ꉯ��ɦ8��$*;&�Sl�`�gc������"F��h�t;��摤�@I8�T����|���U�Ԫ� J[�I4��b�(�m����fu��n�ѕ?T���?P0�;�R��gP@�������b�d�{�m>���`���F��}=�Ə2;C��U�.�%���hf
�l�\��xg!��jR�ʹg��ǰ���%,�Y[ٍ�w&�q���Q���dd97�ѿ�z��ctm�կ��5�/>tH�?h��6d���m�(�LƃX/��2*bM��>�@����#��4��>,��>gc�-�j'$��s9޽��%��K�H~B��e�J��]R�L$P�53絿�Od,w��*�õ1���N!����$���o��$f�~��$�0��WEQ�i�o5X�)�fUP�٥*TM��V�8bF2�+���,ybb!F��`#�h)C���"�|���O�xڽ��D]�i�x*Şu�K'��'o֐��>�=��/�N�yy3����Gq��#�uyHu��^�K�ч��/�c����L_k.\wwS����R�GC�@ܡn��+5���;�Y���O�%U��}3V?����_����������͎��o�S�z���NMx���ڋ/���&rf�ܭXb� :�5��
'��1mD��-�˾(� s���p�	269oיɍS��s����#B�#��oHQ9���2���!`��?4�9�{�Z��RvZ� � ��F�R �"�2mSv.��`�.K����G#EW��W����k?�z�MΦ�����
�H''�&�!Z������6 �Y%�B��w���<'�ѝ&S�q�,?�[u�@3ر��VB�F��I.�^�ўޅ�5]i,<��D�ҭ�@�J�Kti����DI�d���J�B���������g����3��ı���Bi�`�/E��Ǧs4�ަ���͜a6E����s@j��otU�Qq`��lǦ��s�|���M{X����P�@xd0�!dwSx,,4[��^����@�*}���}��Z�1]5��1}���d(�D>��<��:V�`��m��>�x�FWk*x��Zl��m8���<������
&R_B�;�5|,\���*'��*yw��U}^�0y>u�f4��2ː+��/�Rx�,���\He��jѓnw��ߵ�����z�e{��	vޫ��3͜������n�mO$�lŌ��S�.���G�O���}���s���$�з�n��l��j��!��'�yf�t�s���|�<�8U�����z0� y��'�dj�~"��Dd*(?>��#�����ťBbGM�*x�&#i�`��|g���x�tS]�l�s��Xiqބ�2���+� !;[�%�@�;Ʃ��I��!��i���d5: �q6<JC�&�DB(�$�0��/w+�����ǆ �I\�s����O1ԗ r1�Z���$a�_��`��i�$�h����\��J0.?��λ�