XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��q�tRu����D�m� �H�S�[�̐�RF�[�t�h\F�rtC��7	ZV��h��Ab�
vq�JT���Ś�
Z}����AgZa3Q�P���<�SQ=Q	�u�"���|,�*C=_l�[e�y$�GTK+�ӹ�H����>��Z�}�[����x�N��P#��߂����s�F�E��-F�SpN
C�A/l����Qa��W�Y��w��%�t��B����A!g���o�f1�T�C�Z��nG�/FM9���҄:<�/X���� 9#qh�du��ޔ; R�	z%ZC��v�`�=u;�l7>�Qa>���65i4}w�/|�q��Sg��H���e\{"2�Dm��,�WX
����y�z����Kq[� �ª��`�Lv�K\�4��P)��H��P%�N!�÷�|┒��Y7����Te�����@�?�v�Tx?E���+�1lq� �PF�&�=�/��]�#�a�
^�>��>=����\3���X^���c;D�awF���a8�gkv�%�31��RҠ^#$�x C�`��75�F�/�Dp�;|r��T�����nX�|�"�hlȃ��Nـ�A�������l��
�Pi��piKЬdi��4Ep�s [���9"\�!����'8�9�2�-i�ʹ[XC�?U��&�97����&E�Z�����l��S������M������T{�y�A���ަ�������fH_6P��z�2V�=�N/����Mh��w|s6�z���)��mXlxVHYEB    63ec    17e0�Bl��Vk2~GVЖ�=V~�L׷�G���2�F���8�j��\��X�H/Ą"S4���z]��>ȕPB��u4;��7�:1�� ��	,Sh�$�?a�
S�T�h��%T3�	�w���y�ת�.�a�F�z���VC��f�M�V\�����[���߀�dr6��q&�'	`����b� �' =ϱ-	<R��K}*KQ�ԈSv��C���ϴ�_�3��4�̝����]�E9� g� KAK��}#�~��ۏ\��*mB�p"�e(�ElC�ɅlnGC h'J���T���"��]��X����k�j�#���Sߐv���"z�����ۀ�Ȑ���Dkh���ߠX�-KZ[��-���T�s�Tr�?n��Gylx����h���]�O�D巡X	���V~�օ�j$�R���"��K�-%iO>�1�{�"�`�� b�az<�eEۃ����7��jWz��YE� '�AI�uR�S1,��c�-P�=�9,���[���������=5�lS�[uig����C�t^�hϰt�0��5�Wìd2�~Z��n+J.cY�A��8��A웳��g����mWx�9B��N��[іL��#!��v0�<
���֘P��Mqc�>}��t#�)�e��z�j�5��(�|�4f;����E�H��y�I��7�۝4�it첤�*�����q����p�����7m���ZN�/K�o�۪}u�*�de�4��)HI��M1Q�Y*u��|��|�d�I�De�Bb3.�D@���"���'��L�uJKLdk����K��{?�з��@�Q�:_��h֊�d�#�\�(I�5�PFi�weK����U�g�y�?���F��_z���u!�����օ����3W;��(���ׅ��x����*>U�袌�W�����E֟M���TT䃫C6���k`����wס r|�<�&0�U�"��0�2��9D�~��s<�s�A�hPyM47*�;����lP;䮋��p�e�=T�rG2T��[���
�֣�l�paZ�����q3�Q�o>x���%�(�"��q1)��c׭+) +,�OdI8u�c�3�p���&�e���ߔ<b3:��v���3��!_DX�ң����WO{�o�U�VcJZ�%��t�B���2�ɲIe�s]q*�S�n��r�]�]�ܟ�Q�G�9����XT;pbS�K\Hّ���*��Q�z%\�~Q�R��J�و�)���O�#�[4@9U�;��"�,���h?�tp����P+�Te"�GnL1�9#��O�6 Nl�2a��ܼ4�%�*��埣��֌4{����������Я��IENEX,$*�E:�����	�+Ä#�!�Bp��/��Es���PJo�Z���L^N�<R6כּ�z��C\��m���~��L��-'[L}��4[�˵U����۵� ���m���[}Z"f�7��g5�F#��F6�N�ܽ�_P��(�$Y�<�a���G.�ygk����|�K��5"�T0�]��k���Aj-�z1f�/�o�R���c�8v��wz�)ZL6L��	�4%��pL����>�	���
���"��%�]���ن��2��	V�ɴ�&�f����
=�����~ͼ$���j1�\Ƕ��1�s-H\��Q��K�;wPL�Ŧ0�g,'�<����z���Ed��1������6WT[��q�C,���[���pL�+�����B-a��-�d.���X�Al��\�;>�c�j�;��햛*OoK�VM��Q�\�j��Ԭ�d�Ϲ��ӍF��7�e�B�(�@����|�>��ʂ��y�Mp�\2k� h=���;��u�=sw�r����"��V5��`)[j�`� �=����Q�lmoH3�Š)�On�L�^�V���lǲP.)�_��y#�r�|"1��m�J��b�
��}	�
b����~�iT�c�(�8(����-4�Y)�M
p�K�_r������[w���t�Jƹ0���+�u�-��w}�29�����=�s���wd��j�o/U��0���` �~4��V2=!���-21�Z��8��-~�3���3��t��ն�*_�=�=^C�V��!�1�͆<� �۔R�]�
.�Y�?7R]����vE�1��v�6���|����T�|��>E� ��y���\�`�*���G�@~6�[[��2��бp�zF#W?S��&39d��\�*��~��b� ~Ʈ�~>�PGI]�� �-�eh�"7�� �e�g����Xg3%m����A�k�H�A	���4v�D�=�^�=�%�9X�mv��=�2RI}򫴏��^`�T�]�Ze6��?^�]���s5N��K%U��E(�~�G�]K���i�'�ۛϽ�>�\$}т��`[[U������{�� �c�֥�(q���Yp1�����acX���>�1[�)�E��H�GD�8Ώ�~,@Bf���u_�W�Ϳ�!�ːFH��s�0�A(��O�H�t�FT*�1��@�׷�%]aǲ�5�r�
�K �dj��4|ֿ���͹Q�\�F:W�|�����0;�\E�`:[��{j���$I��N��=�Ȯ$���=M�������|�W��Z����7��t
��G�l� �4���y&U%K�r�� ��r�{���!y����5�� K�q���#S�s�� qd�
[Gc<��B�������l�x��F�mfH���6\�p�7zŭ��d`f�ٜ�����)���(��� �M�M%�m�MbcR�{f�}��<�u�RΥ|^�]�? `\��?q��+PL�~�5O	:f7z���2��+SLnJ��Iw!la�g���c�8a�LX�H>��2;�+BP�/C��D��	$I�_���Ϡ��NA���SU�UgX��8�B�*���{v���y.�J5E�LF�Ğow��h5D���B���ԌQ��9���N�y\'zN�
� Xǫf:�l�'�{L>��sYj�uǡ~������\B�Uh��Ҝ_a����S�)	�mj�"��6Wh��F�~�g�d�����kl�d����1��@���'�Ml��)�3Cm�	�E��|��T��O�B'g���Z&��Y�6�O�������@���b��m��g�D� B`�C���H}j���r|y�c&���h�ɝ�!�l}J��9NY�����(Gǁ�%M�QwM���QF�*�p[L}�~"��b�w� �
6g~��؝�Ӄ;k'�=�dr+@�lu;�s�bF��
e"A��ЯV�&f�c��=��5}"n���w��	��ԛ���M��Lt��>��5�A5�3ce�cF	ͤN,��}d i�i���[+���sI�֑cA�6ob��s�aii�ȿ�m�vC���#ۜ���bR�����C�# ���,�*� }CЏ�?5�K"�$��.pC�T�	�����oE�K �j���5�-��T���7�A£�3���0��"�:�Nc.ڢū��f�#�ˆke`�u8.Ǒ��m�Y��8��	�	��ءo�t0�������|N�aˍb�����K/<r�7X'�U"�Èy�����~�	P(��59�X�����d�=�O�>�j�c��cF�)'�e���֕kG���ʭ�_ӡ��k7��b �bC�n�? �ߊقc�;�Y�.�*�81���w@L;�^������e�z�Ci�!�3r�<P�03k0���8�S���S�a�2k�������%��
j��GC��o{_J��NO?5��d1�#���e9���'S,<ɣ�R�m�o�h���M�Fj��aP�E$��M����l�Z�l�9E��&�?�)4�YS��,��>�E9������ð�\���"�[�?�^@O�:���w�M�D�6���M�u� /-���g����;5��5ʙ��*x 3��x]KL�Zd��BZ:(��Fm�C+���U��� ���2�(�[�y[y��p���!Qn�G�'�)9�Ń�>�����+TvC�̪�b��U�.̌�p��:_��bS15qZ�����~��hn8��k0Y�g�R�4����1�	�tߊ�Ȕ�i�}�U�^�X`�jG����bM[s��dA�����̙5g�\��=�md>Q�<������(7�ӭ��a��d|6�F� !:( xB"s�j��������[�m1�^���.3dA/�:^�d��Q@��T��Z����'~ˠ$�)���y����֍-J�KD���p(��������ʲGݸ|
�"d���}ԟf%�1���Ō�R��d\+�J��N��^qȄ�'�W��K�S��O�h�\�^s+�&����o��P�GM�0��xL��2���'���q�)ƌ7����x#��`�;f s	�f��n1�u��О���z��K<v�|N���x���yt}�3C��T�Ckn�R��S4�6Sݳ���?ux�f�*���Qo�NR����;�θ  6�Ĭ�#'��V'l�l���`� ��7�9�-��p3�#��|;��omxA�ğv��sK�`AMq�L���b~T=�`'c�gD�;�>���Za�i��i�)N  �Ě�U*���e����<1�K�.�q4�"��Ո�0����]�� ݯ��J�y.!P[��q���}{v�zL��A�n���l��<H
�׹@�h }-Uue6L��/��c�|'д�(E�1��n|I�&�փ���J��З����,te�!A,]�cڢ�Q��[��C^IY�wa�a�I.o�������^'M�jфE�	�wT�?�4&Y�c8���yRQ:�L��� �O�Ѣr���ܦ��G�Pv.F�U�y�4*����c���v�5\�on�bɱ#�p�TvGV��ǱG�D���x|�<�Fk�u����H˥UX�(�3�VU,1_�F>z�����q����2s��[	j.����6����A:�Ј+lEb� ��h0uO9�����-k=�;Ф�]�{���͠+��m�lM������q��9~l��1��m�袰l��q�����q1��}k�GҔڿ�rcP�^H� ���N�_�^��J����+(�C�l{�)[�n�6L#���D�1�w�&�0�.����h���q-���n��0
�w�Oqӊ��SRi�'A�1cu�i(l���A��������NMQ!���g��E(`ml�jZ����Î�w��'�j��_�@.�P��7D��p:���![ㆱ�6���~�,�೙�J��)+�e��x�0T!��{\tn�a4ˤ�/�Uu�����]k�P_$6$�*��)�ã�E:0��j̵���qQ��T�v-
�?g�ON<a���`O�`����=�#C�!)L�7�o�b�bI���%����s-L�q{��i�(� E����*�nh�'��&n*����U��������a�G�m<h����Z���j8!!��E6�3ǹ�}���"dC���/g�I�`Ǡ0��4N�;,�;�j��I#n�������t��y���n���>/a�1�~b��a�Q��E������#�F����
�?���
\5ma��mS��Tت%*�K�H�Ƴ(�=;	���OQ�B1���V�w�5MZ�T�_A���Is�U
���xͺ�S�<��p��ۊ9f"s���ޣ��q4�K7�9�0�aW?s��)�C���x�26�{����١���%e�yMy�d]	��.J�z��Ʈfq�\X�������ʌi�
��^>#�gU��B-�����k�[A̗�h����љD/�^*h��>$/=���9�V߿�����z9����5�F�PO���\?�PH�U����)�����Az����<L]$� Mmu�T�cq���4�mDq���xF�L����� �A^����kL��ʔ$Z����q�Im_�l�胒�W�ʻ7 �1:��8��;_H����3��Lf\��ֆ�