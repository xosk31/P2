XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����SȎ;��V��%�B�&
kv��r�Mg�W�7�M4u��NՖ$��^y�c�����K?Ջ ���z �'��S5g��u�6'�
��\�u����O�ӡ�{����n�6n��*�8��0���z�D���RzQ/�<�8rփ�O�N+_�H	%G�%�I>4�O�)Ӻ���~�u�6�%��!亱�WG����~�S<���vd㎈��N���J[Ⱥ$ֱ�w��Ȏ�G'0:3��#� ���oU�AR���f׺]�e �D�L�J��z	C5ь���2x�� �Qg�2@�u�W[œ�w��?2��'!�Dep>,V�#Oh�ю�x2-8���[ӆp�s�dn��I�/��G��gt�c�fj��n�ɉ~�<¼�чo#ك�?%��Aڶ"�J�+�Gw�j6���q��lb�Xs��6��c|�鏻���2gi7�/iE�Pes�<#��V���"oΡ�V<T�b���/"j-�Y]5l��Hv5���oPA�RPmŻ���E 2�b�3��
I0�/����DA��~���"&5�hf`��fH�[�:z^��el�&#��7�9�/�ÿú>�M)di;���5y�hIԴv������� ��̘�!�RV>:r��[a�x�a�m\p�u���ǟF)�پ8E��æ|�����k :�����R`��@i��lU�}��W}Y��g���+�jn���������xΖ�`쇝�@Im�_ڀ���m�LS�QJĂ��(��q��?�r�@��
T�����s0XlxVHYEB    fa00    28c0c�M �n���^�\/N�1Ldz�^2D�J7P&��s@��Ԣ�|�0Y)���/����8��
���.�ll�{6�H��S1
�)����˹X��� ��>O����כ�X�*UY\�qh!�b3`SՏᚆ�"X��С\�A0c�`�9.,���۲�M��&1v���eG��-]�L�M���Q�-F9��f����4��.�D�1IK��'�)^&�el�,��7���M%Jrkƨ�ӷ��T?f��5�](���۞U.���2#�^k�U1W���	vJ{�y������o�n�'e�܅��2�ە�����\�Ԙf���D
ͺXG���18���ݖ*��t�"�^|Y�迟���>��"K����Ώ���Ŷ'�^���Wx��;A+���c��،:��^��%E�z�T)H������+]�k�S�e�?���j�2����۰n�4���כf��-$L�Y:4�/u�N���P��W�p�f����+�|f6K�0�����������>U�@�h���A�,q-劰t!��o��S��0��Y�FԨ���ǆy�+��6��C��q��W 9��'�7�;�o��z�vD�]��s;7����fv$�|�q��C5�c�G 	4���/�k��.��c½���r,��Y�9��7
X�5����OW4�� ;���<ը��7��Ǐ Sr�S�A#�Y;I��20�%)O�o@2-v�r|�LU&s�hs�}>:�]�I
�SYQ�Q�]�6~���� �����G-7��>'�ӈ��̜;Z%��㌛�NY��9	��� ���]�ԞX�NNo�)O��� Q�N���[ɥ�?���?�>4����;y�2/��x2��T70i�q'�69R���:\ ~���x�AP/�O�~������Tv]�({���*��zL��%��z�/1���J(u-|�Pu��*��(z�x/�{��9�U�E�(��R3��*}����n�.-߯_�A��W�	NøIG��|�l�l�Jb[q&�iL���� Q�n��qw]�B
P�ϭ);s7��[@� �%��r�ܬ�J"�QO�L*��<�hQ��{��lEH��B	��|��������C��eWo�6����6�ؠ�����$�.�~��"4�U�}nN���X%�+\D����Xw���zw���M�mw������\O��dU�q�����U0Ϥisq8�5�}�lUvo�A�R9=�9T�����}G�Q� �N�^�;�x��!��^�ي��`X����d(����	*�P$�F'�Q����a�)\u�bu5�	]r�(I%�������/��S���a@Ha���ǥj�d�0�ɽT"�U�(�����Dwko��-��&�K�Zӯ�`˽JP����Y�b����2^�E���t����C�:���g�i��-
^��w���" 5T�_�_�	��Zxɓ�����;R��4h�Wυ@�r�����:Ѻ��-�o6��@d��	ކ:��'��Ht֓�JF\M�xli6�됋n�A����H�mDV@�3�m֧b2vPuI�����\�業���~;z� �Yg�7ұ|C�,5Q�OYu�\�������ї�ծ|��Zh�M�v]����PB*[�Z��ZԆ��>�9:R%���Wz]���R��,�N摭��uڃ፮�~�ְM���ݚ���"�2ؽ�e}GwM#E�'��.5PkxřF�z�y����8���s�#�s)�XzO�$����W�5�@b����y�j��kv�:��0]b\_�pK��bw��6&�v���S���&�#��&��J]�c�6��l
}r�'�ˣS��@�3�/@`�ݮ筅jF]�D��Ӗ��=�����`~r
��:h5�g2���*w�lD��2�@)"�f-@r������l�4�/:�A`��l:���� 2'��Gqv_��o7�|�[ ������m4��)s(��_Q�t�*�
���p��~���\�_p)���c�z̶c�a�,@'Q1+�f��}�S��^9e�\]XJ���~��r���/�	t���zނѴXr��Hu�8|��.\Ut�A�D�0���n��#�T;�H�~}~�5�U��vmi!j�o"
Y��v�����Vj�oOz^�@G=]{g�]z��R��<��Ll�%�M��Ǭ=7I�}xQ@����D�� �Xo�K��U��WV�}Gi~i�/�e�Rk�XE~Q��)�����+K�MJUAm�� �\�4��hzS��
��@��-�b�?�]� c$Bv ��9�<E��z�$�c�*����(:A���>����PҐy|D퐙�/q��-��vw��c�>=���sm�O���6Gu� �}u7l�LwS��!xKx��Ɋ&�su,�OJ4�A�n�8��׌1Xn�AK��C�0#r������U7hwr*;>A������hj.`�7	G��GTG�RP)�,n��C����`4���BӲ5H5dAŴ�s"�.�"�j@�jR���$.Y�ۄ�Z7Y ��9�`1<m�	a�͋ �/�*T��p���}B���v�,���a�<k�׈���%;[2Tzma5��?�b��;�U:$w��;�M�����-����5j��M��U��0�av����'�	�3~�O/9�̫zk�{ǝ~y�B�]�cU�Pjɛ����V�>�� baZ��CP��~O��Xi�u}��"v|P�`᪽�q>N9[Z� £�I��l���,q)o�>����y�l`�Sg)�^ܔ;��s��|� Ǚ<����m�$f��J���p�1t���L
\��d�#ҧ���D�b� -�ō��H�4%�:�)�����.�(�\��Y,�W�b�xA=v֍�A�۫��7�g���+�͒��hQ�f�Ȉ��ϼ��A�G?�J8I��2ePA�*�w|�����S])��>��_i)$��|����}�S!���5��81����Ǯ$����R,��s�L0�6�sI�s�EŨu�x0�#ZJA�� ��# R�򱮽p>����TR���HfS���y�Г�o�P�JVW�Y�:`Σ3��մ� ���h�k�"^f�x�튪�C�*�-F�pZ�W�~��W@��nL�p�s8��hJZ[�S�G�=Z<7���X M�9�b�,�a�򕲍XS_��~<���[�VY�Syg'����>��	��4�6�m�v��H��pxsk*{h�M/��|�>os�߬��XXA�.�_����TYC�]��C��ZN���.4��wn��Eȯ"����D�Ԯ����;��C��6��`���+5�;��Zn�w$�ۇ������v^l��zF���5����Q��/;s�Z{�̜��p�Oưk�m�̤!c�t�}����!H6��<�t��Y�ϒ=F��Ww�,��i�,��T5�6=���3�M5� ��|�����\�b~A�������`'�u~���U�p�`�%���t�~,d��ϋ*M�1rVcO(U�M�w�(�"�
��5?�����k�nm�R��_�|}�i��g��O@����N���z�g�$�Qe�24	=��+��C�el���;��J�"����(+��E�Y��I�gpV9�<eSB���t��F��~�ٞ.����QR�3n��jH���j K�+�mP���M�6�G�p�?�4�]�)pӗ5r��I��ͭ�V!$�S2�d��3C�Y 4q�ߓ9	��Q6���.�m�a������S�	��3�R�	�e��b�26��y�$����>� ����t�I'��e$ׯ��{T�|�����ǹ�WZ��� �֌������_"�F�#TA_eo+���H2M�'w���i�@�kV�z�)�?��xha��?�yA�QD�vQ������JYRSH�Š���e����"�E�}
�1Q�M�xl���
kx���O��_U�XY��ʳxb/%:����J����}K���I7�i��Ψc��S�׻)©'K3M���Fj۝240G����H~Ȯ��~g�?�=7����K�%(���=���'o&0r,�a#�A'��l�@��-߼���W6`V�!�� ߭���SB%�Y���k�2��󼮵�Ï�/5e�w��Ij�6�B-WG(I���dg�K��3���%)]���`�ab���m]�ʆNy���K��?��)d�^����w����@u���.ǲ��5X���KϺ2�����%-� 
��$��<�{��4Y���jW�*�mf�&�E��z�6jȤtC�r��9������@�`�wE���{I�1Y~�DL�C`���w���]&����2>�+��^��mb��jЇ:��{�@�lq�͎
?_�x�l8�聠�IK�w�\�_������rJ���/xs���NWAQ����٦W��9�bNC�g�.f6�뿒���;q��>�~�ʲp~���L'��z�d�1K�ݯ���\���g�T����ƥ��+���!vads�!6-��3b��BsfБ\gNY��D�`�]u�k<<�I��̗�iʸ�7��L������ܫ�|2z)�@*ω��4)�P����	�5
�9��!�].F�T��Tg Cp�I���H%������f�h��
PՁ ����HR؋K�ܒ&���c)qӯ��Q�3�F�Pj��1ل
�ni�H��i�ϱؑ�z�}�9��0�1c�z�T��)�ʈ$N-��?'c�e/���k�qnQ?�*l�1�V�7��U��oz�|��c5�qf*�T^�
���Ƣ�P5E�7_o(�*�F�����S��9u������K 8�"z�^�:�����v,���@xU�^�YH	�i�K�٢d��x�3Ȝ��� ǆ7f�$q�B	m��v�۷A�����X�IT�Y����D����?�G�l��J+3���Q�׼.�lA9'z�M�^>��+�0?>_Et��2{�v����+A[Sѐ=\���F�s�����0���d..0+��>�����~P\��8$�Ԋ��v!GT�K��C,����i�����{�W�p��~�em.����uYA�󔣩`N���v�BE�hT3hň@�<&�T�'�D�2��h�D2��flQ̚��s� V���r}&E=R�ܜ�V��������b����󍬫;�r�}��[���2�f��"s�J�)V���{���T�v>&zw�]���0�I��&�W�=�0+���&��H��H��'-$6G�ѵ(uVQM����}�6ە�s��%��9��%Y��XX	����ڣ���m����Ј�R��t5LI�=X�.)�n��f5�'�&�_���j~cm"��+2+�H�)9�����8\<�<n�����X4��P_PM�%�-/�%-��ܱ�."�2���`}�U�E���n}�����\�iɒ�d�OϠ+���C������C2��r6��?���;����f�@�_�s��.b�����/�����������/��~�i��L<�7��{T0�D3����	��È�������~`5���%a�l?��Մ��t�]Y�����o����i���G Y@�f�[b���� �}ζ��ASEkrq4�F@E�p�{b��$�2x"EN|I ��~���r��08l4�\Yj潰� ���������'͗b6�N�}��	4��3��E�dk%+�d���Z�����$�w�ւ�Rd��>5Q�Y�^l�k��,��l9�<���]WJ	<��#^@�h�X��@ř��q��ª�=�A�{����D76G(ԅ:�|�*�2���f��B���u`�I����¶�'t[5�> �?�� ��L�A��|BL�{L��Ub�J��o�Ƨq3n!�#��}��)��5�k`�s����jE�`js� NK��M��č͠����9��N+�$�����[~��4�`9H5���s�-u�K^v�R�g�D�"K��(y`߃�w���[��Y��u(q���Y���Y;���uur8��@rj4���X��U:$:\1��m����꿾���u�s�]��5G Њ���[�MR *�����O���`����<��l��D��4�˹��B�,�t3 ԯh/��?<���
j�|ѻ����=5���!C��[�!���������S��
Wf�E)�1I����[f�G����� �c)d�u\J��"�kϴk_�b��ʐ��!;��?���6�0��⽠��-�ϋ$�%ɜ �f�V0�� "<��c=ZhO{�?��88��>�i��[Y��m�V�XN��G�M�Ѕ�@Fj�7��� �w�IJ}?{(�!Y`"f�{q����F@��0Y��~�#����4�&Y5�.��f��ߑ�ɋ��ߪ|o�e����X�YQ�s��E) xO��`/�]���RG��`�9K=i��ř��u�+�=�=�"Ue�V�6$�ĺ]vrm�NS	Tl4r��0B�g<�ip|3��d��A�YbT�л�����|�&��@�m<(v�;f�D.pE��R܏"GJ
U\bu'!?;{Ҡ��ט)�]�BB����Z9Y�Ȍ�U��J�i�d�O�t��'�� ��m�v�B����*��]�v�z�җ��'C�a1��.�Y-�z�R����nS�p���7	!e�;��`�Y�
� �Y//��M� ''�Xm�$/�F���=�/L�+�v2���{K��sm���
�d�����@
�u�&�B���Y՗G,��\����j�x�����	���[o_1�� �r�g��͠�A^V=b�E1n��I��4 ��Wbo�C�Tۤ�nA7;*�U$�k��B
����V���N��(����T�7���)��ŧuHd�AKmZ��+��8K�2�O)I�����o)��M��(��J�d����XN[Z艼�i��ɓM즲����������9S��O�@{\��y������q0 ��c�?�s���!���ʖ�df�����km+F95�ט�>6R��bz��H���r�z����p�����.X�nd a�p���Q�e@ѧ)-kMs�R�6�#[�f�� �#�\N�&*}���s5_���� C^��<�F�����\�%euj6,�t�[Ծ��@ԋ�k!��2�����Zτ��>��~�ȿ,���b�^�#D�R������C�/�%:�7�E��b��ea9FINB2*Z:�����: ��8�u^x�Ќ2#�s.ŕʢ��S���H�$J�z��~�����޵�4L(��Bh8�ZP���ʎ�$?X��5R�,�����"�h��$2�7h��r��-�f��S��"�Kl�n��r�>��m" s�	���a*����qu�k�(:!e���t6N���֮��z>�55���{3O��T@�y�G�s�셬��Ki��H_~'Z�Ǹ[� |��+���-`����+rf�I�n�9�����|����-5�O��r��'����sɌ��%qS\��c�uK��Z�����-U�xAf�
��ו� c�����Jlp�8�F�����\뗯�1�*]m%�jm:�Y�ZM-�0޲����_]-�����C1x^���dꗰ�B��6��x
o$�]a뚪�Č�~��G}�_�:,�1�w\�s!D��l��.5N����
�<o����n졠.4m�B��Z+�?��{mŪ��1ԅ�kܷL͉���XY~nv�	Qv�L�b��L��qu")1��4f��.EX8�����@�d�Bv��C���H�.�Lp��,��Ss���	�5};íX51���WL�w2�/^Bs��L�% E�'��6Έ�U.w@��z�ϊR�>��K�B��r��	�e\�W��\>#�V�X�k���~C#0��%L��s"��H�I.��J�aw	�6����U�=���ir���6�!?�<A��O]�� ɣH����{v�j����(�cH�9� ؿ�ޙ�K�+�H780�����5q#���X1�����S�p(�R�����X(7v�����40ZVS�q�6��#��~�"�7�K�b���E�[M��1+$~����T"��4�ڏm��Xr���������=&}È�u����(z���F=E���Eyޓl�,gA^�g��(�u��Z�3�5���q��]-�N��r����pa���<4�̅��R�����ǃ �KΎS�=�Q�z�A䩈���2<Zm�͘�͔���K#�����p�(����Z7L�Mڝ ���)S��}C��˷,3�#Ŕ
��3Y��[�T7�:@!���#x�K�
7�"r�v(_�-4������*�1�.�����t޶`���`�	�xrEq���2��XU8:�uMqҶ���韒��+�õ��1%9�+��2�l�	c75��b-�66C�m@���,nåA1�R�VQqM|��n���U$�q/4{#	qƦ0Y���ӽK3Q>�$֗#<�Y	F�U�ib�f�r������S�T���f��F����%Wi�!ԟ��5�����Pg�0T�E�l䯕����70kT����'�O���D�5MɒebG�HFk�����~�J��Цݽ7O�>�����n��JeH�)�'�岙ʖ�,Yh���t+wy#3�,.:-�=$��s�A��X6%���U�N8���Y�M�MȀ���4BG[`��ǁ�a������H�*kY�
o�Dl3�w������*�&�� mi���k����L�X:ֺz�ͳ�YF�˵����$�����V�g57�J���hR�P8�}5O3���&
�x�Gd�p�O�Mƍ�&?@����BWOpt��T���`F�D��G�AvY̆{~Bm����o��)-�ŔR@����
�Ν>�f--���C��������1 ��~L
�@i�|>����H�<�H5^�esi_���K7V��"�`��$�nz�u�h�������h���բ���"�>z� f�;�.
�,�B4�� j�d��?��Iw,��Tȇ`t����kI	U��Mu/d.�#�ʣ����(O.�c��(����K5At�۝?]=|a_sQ�<o��K!S@�x[Jb�nTж;_&�d��6���3�|���.��'�qsm�@��!^)������*����ƀ7A[�/s`�[-��l-����>>��{*֏a֒�߿
hL�c<��eOy���<Č�e@�R���Wk0�
�-���4a���j�~&&��.�\u蛧�����x�d�����`��a����P���6�y8��ҝ?����"���I?lSk�M�ht��k��CV��-�M�����ĉ0���I��S����+�`
_De<�#�zM�i�[_�UD~���4u�x�����2���j^�Fi�0�y��ҿv�#=�E�(�mx���Z�x�H`F�&XE��ڑT;���Y�َ�:�uwEq?9�qn�^Ik��M�^�V����S�S���"ϊ�w�?	�~�06˲��M���q�J��9��M��°�JMS5����15�y�jd�=z��<-�^�1b�K}�o�����e|��y�KD�[��dd�ozD�l\$�b}Av�v���$� �#��_��NsA�q������B8E6���}���u C�;�� R��`�$�Q4ѓB����noϙX�����u
�*x�rݽdv�"��l^��)�����],��!fYJ���h�lkfJZۃ��k��
��r`�F�u?½�T���p3:�Y�ɺ�A���Q�o�'� 'jR]n7ϺG+�`��'c)��0QS��ݸHf�F�ay߻���[�4�轔p���I.��4<l�Է҆�n��c������68�rL�;��lp���<�OНi�֝��k}]�����];SIA~c��8DC�sT�8�	N�li�P����ڹ�i�{��������g�)F�i��[�e����2�n����8Ŵ�F}M�=u��5�Yc9�{m��;����r/�ea�ەP��W
�I- �[
��6�ʤ�F��-s\����uF+�˯��z@�����Q����oߒ�k������Ļ.�>�/r�=@9�
�r#XQ��X��(�Kl���OY�������~|�2~��p���u��Ъ߽��|��u�Z�&.F��!Ƞ�S�'��p��+�]n�Aa�X�h{�E"Ղ�
T<�p��,x��er�&�4����=�-�voD|IZz�N���Y2s9�ٌ���a���El�N9��<����/p����P#<+�,x="�����j��1P�p���4�SAQ�"�q���ȔI�_��XlxVHYEB     896     280�:Qt�ZfF��M���eS!�m����@�+��zn�q�NN����"�b��:V�"�X�
�M	{�̏Fkk�gL���	��=B�Tj*s�ҷlU���8�V�"[t?����{j����p"�l>s;��{���\-8���ňt���k��.��CO��qQ>O�r5+s�8�&��t0�ݟ��q��ؗ�~�ɿ�g���4g�_A�J���9�`Ė�.ex�C����Z�IF&@�};�� Hc�¦
�N�fo�W�c�Cy�Mi�<����s$���ȓj��p�ᆦ���J8���o/n�*�\svk����>�ߥ?���Q���f'�s�����3��{.֣Եz5��[�⏾�C/4�� �F�4ű���;�׏�C
	Kȭ�E�x#*S��@�-@U�I�	Z�����K�)a��s������+`#I2cő�<�v��������������w�NhSA�Q!��޿-qPb�A�R;����>A�3E�b{�4�Ǚ�Q��h�\�������ǜ���A��҂~N�s��a!�����':�|4U�H� 3VD�]���4��vr	���H]l[�ג�4FI_�_�
��)R�x����%n�^��d�>�d%l�;T�'[
��