XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��6�"3ꘚ��M��GU��C��&]�d� �7���l�e��t��P�g@���Fە5�,�YJ�U��-����"ʨ�hx��Z���|�%yj���4w�����i3N�O���!���?}X�M���P�k�M;���	�zs���f�Qc���S��<[�yy�%�}����=o���f�C|�����\��N�.ˉ�UO�L�;+$���D�H?��K��Z)� GΡ"��qց�^�#u���6�
S�����z"�
��@�Eja~Yߡ<	��6==���Z>�J[�ߢ�R^��5A�V����T��k���CC��=���"��x��F��U��/[4��)�!��d��EMe*�E�� JK[f���}-�v�oI'S��X��+��H!ȊcU�T���³\nQ�*i��(Ȱ���	��_�H}t���S�d<5�ϖW���M!�	�R�鏇<������a����sH�>U��6R�+������sP�P����I��*�A|	����q��;36�z]67�ϝ��۩ԧ);"�����UQ(s�eU�
5	�,4���~T��t��e���}����4�Iv�܍ �\�U�]�(ci��>Ӑ����3뿊K�7E�۔�tȫT�4�񉵏+����ZLi�Y��F�
�<���qx��*9s���^�C�Thn�.�W�˲~d�O��nB�7.�ɪF=���Qg�4�7��d��-�O���)��q��m���01I����Cm���ޮ�g~Mc(XlxVHYEB    3099     c40���ˀ+�K��Xy6i�_R�Og�w
KY��~1j�b~��OC��n���V��Y0)���?k����x �Q��Wd*y��hE#��t�W�Y�+@�}�JAX����tے[�\h���+�ik�֠���:I
�	~'k����y��,ē)��xX�Ȝ=Gb��}�����|i����Zz2ΜB���M�_�5,*I>����3��Kz5d����Z�?�p#3;��t��PO�T���&L�L��	Èp��uH�����h�\=��0n�)����P�,�\�w>Q�����_�e��	�ʚ���F��a�g���#h�R�I�{9��!��v*a}�)\AP��(����o�.��V�k�EHU��h��-}�QGL�\y�}��&�5��V�A�+�E�i($r�!���GkQ]`�Ѹ�r3���M�$_M�6n���j-N�n��Qe��kxsY�q���e��}�F�K��𨂬��9e�����A5U����I��Т�F��\�5� ��e�m4Q6�cI�L�H ���A�d� է�e���c���|��a�� �t��Y��I��Ae���w�-�h��dC�pbZHߍ#��Y��֐v%�I���R0�����
�'*�d̬��~���6 ���죌�E\���=��F[�$�sd��bey\t�㑈�W��u'b"��@�ǐ�'�Ђ@M��Y��*�[��Opp���s�B��X��"�J9$��~A6��]t�e�h裗�to��<�φ� �t��[���2�d�}�l�^��s�?���݈.t��ڴ,���"�N�M��V��
�܅)�����D����:���ڴ��h���ZM�����K�&�R�LJ�$��xSPD� ��r
+
[n��{<�o�{�FpE�+��d1�
"��A��؊/#C��#�M������~kH@���Ģ��0#c�Q-�s
^J.X���� LH���烄-g1 g�"J%������W&���������&S�L��M����T�凑�����)����4�nBוM��p���z�M�b5s�K���p>����a��K��7jw� ߬�^�B'�������AU�p�ǮR/	ľ�o�N�h�O�qb3X��n�Y������)Wno�PAIYG���!��:L�9�X&� �GB�m���v@�rT
m���%��╆���	��n�|2�]p�v_ Y���nHqk[8��� ��clI�߇kZK|���P�M$�.hG^T\O0�A�f�na��,
���s�
+�_���;`�j\�# ĸ�B�	[��nߵ�(ٓ����5	5&�(n�I�E�}k���wuO�܂���?�A%L�&�4r������z=+�/�-�1*���o�;P�!,1)��t3m��9�[��#�x�8^b(i20%����������l�2��i��;�G(�h:�?M". ����D�~Gǣ��ك����VW=ߐ� �-�f��"j��8�y�@�µ�R�w1s�7�m�/�4n�Y��r��/(>U�ɭ���e��	ɜ�"����$U�V�BT�|��Q�4��5R�L#��	��oV�F}%��/�q�ݰ�	7p��~]�H(�ƺ�#}`��M<�����в���M�&�&��e)�r�m�&'�=��9�����ʄ���󔇠�ch��=
�F r҂#Ď%b��QPSD�1zHd�{�c}��=K*���_i��u8*M��zJ^�l��G��ZrGEj*��V�s�<#�؁>��m�* VI���Y�^�$�Ju�B����҈��u�8X͈`ܬ���M����>j���og�Zĭ��8�'Y��ȕz�#�z0t��I@N�|�'���{+���>��i)�ߘ	r!�f�]A@ͥ�Di���h ���H��`�����O+g��i�?scrEI���a���3>�#g��vؒ��4{��ʣ���w/�\|`�q����K~,���b��S<��� 錞]�����f�'� ��YiB�Z.�v���q�?6��ﺗ���h�\�����*�o:��E�џ��,k���[��,o�^��F�<^>�G����y����rTQ�jJTg�����HFYef0UdBݙg)g���X��5]�ᗒ����*c��p6B�XD9U"&�a���%1�u�
��|݀qop]z*9�N���F\���0N������cZ�z��/���..�n7�W�J5��UF�gO�ׅX�`:�Q<	���`�G,홷���i V�d�@1d�v��}ܞ5��o��l+N�����ʮI����?�������k�ӁK��I2"�<vN����R߲��2IE�7g��uНŰ��뙎�3�P�������S�4"���o�Jk�z�h���<q[�ġ�H3/�����,�7��A�̴ /��j+7�Sx�/�G|ĝ����z�&�/]F�t�n|ђ���J9_��a,�E����D�2�B�V�I��]�����S���E\�Rdи6����X���Rl<�V^\Kc�b�oJ��yfP�����0-�o��f��.���Kso����� ��2r7bj��'!æ�s�O�u3��N���G�r�'4���Z:�o������ G~���dR֭���x%���!�އ���������'��im��������Q7����}�n�vp��fR�@��(�A�d�1]��_fiy�	������K@e'�+a��h��E�3¼6�ж���>��C6a�$��B��O�}ЯI��
�G/��NV�:�ۣ�8���xJ2�������+��F�Y����S�� �����֪�A�bwDc��Ω�y�$$LҶG�b�P�j˦%}���๛\0�|����Ԫ�K�~Gt�VJ�p<��4���;��nM+�j���+Vp��WD�����\��V2� �%��-���]��SfΚ�9>[�`����C`6H0)J^,��Y�Tm����������r�~�m��8̺��KžR�>����0P���N><^JޠOZpF�`~ۗ��U/���D/��W9<����|����p������TK��.��B��O}f