XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��6����/�͕"i��u6\��4=SK��� !}�q/<W�]4e���פ�#��|i:����§�<��i��.�p	.���?��jukJ��	)ٷBZ݁%��*�1�{����{�
���7kG��a4
��]��u�s�A�P�@��r��;�޹0#�����${N���WɔR��j�*LI��nR����c�}�ש��\�_���?�ν�c1U�:�3�~KȇTx���53M�<���e���x���<���A1}�ᮯI�Mo	� ���Ί|E��{A[Y�m��@\�����P��-���-~��å`2N�n��Ԇ�p
Ľ'"�d���@hz���:Ro�Ey���DDd�x�2*pn8֡* ��'f�>��ȑ�,B����|�_~'ٶ%=�ϫ�u�L�x��y��,���� [HK�R�q�	���%�>d���]'L�<�;��������|��k�"9��;�1��S�0��~����� 1��Ϳl� 7�dc����Ej�a�U�Bh�"IҚ�ώO(2�vɨO��q���Kxm�Ͽ�r�&����=��¡�r��	�O�ܒ��&�tX�j����RU52�; ��?�e!!��#���`��'sE�eP�?�R��ޯ��E($���+��v�f��Ù��;�x$޲���dls(��Ь�Q/��W9�&sO#;��F�//�WIN1<�����籑n����6�u7�	�g���vJ�p�����zCHj�W��=�m>�XlxVHYEB    1192     750�ǩ(�":�����W/-Nb0�߼�"ǒ{Cm��c�|f^��q��\����<F�����b"���������/�Ad����8��U;%�?���\a������ﾚ�?]��JuTurO��'��
�,񱴱��ѻ�Ţ�kzt_ڮ�uj�y`�'��	7I�\�0��I��^��س�\�#���3�ѨتY�P��O�MP~�=*f�(x����j��x���	��xCŗ�
�����Ex�X�/����К��8���4�q@RX�p�
�6W��H�s��̇X̗C�����>���m�rt5ߩ?􊶣�a.�0����s�G?�7�HAk)-�
�V�V�`���i�OQ���.:�F��X@����,�˟�EP�y:�4�J����y��J�o���c�B?�!�,��}K�Z��Y��}�/�h�y>3���E���CK�s�>Ys�u.�tnP��q��4���s����3�WT�󃾠����PAJ�a�HF<��ǎu ��?�Ò��O7���������H�x^m��,gzj�(�A���]�n�� ���_[��-x@_�{��K��[R�[(�ϘU�akuԫD������N�K��I��k��$q��#��(�iY0�Oq��f-����ؠU��zE>:��~�dZ�t��s-IX4�D��h�|L3��K��I�<�x���2��;�
�s^X�R�4��r�S�S��[��!�폚V.��r��<)�_�,�,��*�Fda��KNb����Ԣ��p�,Y����l2�i�_�0�if)ht�?����e��0L�&�Rv�����)X^�����3:�)rJ�HϿ������8tX?adC@��sr��z�L8(.����G��d쀢 h��߿���(�kě���Zu��V^��r�����a������^v/��[�˩P�}z���w��<�˜�~��XL^��\���%�`��f������5@W��䫶C�#�\FLU�6_��k�8���D7E7���B=���}�]�A2��0�0
�jJ6=1f*Ո���z�_�[q�>~ ��hDf�s*&����q�et��ig?h����C�,�h��qS���.NsL�CY���E�V�r��ʢe�SZ�{O�q���0�{��O� �]�^��ε����v�@�XK�xW @?�@�Xq�TyO@�
/��~����I�/x~-In���a��v��f���!��Z~ \�x�f�,ni��)��"����LI�
��XԬh
��'Ů�t_���y>��0s^p\aR_^ߣg%�[I ��,a�Z�p	)h���h$�tBu���sߦ�TƧ���N��ED���9� �q>��f�`y����n�]\���;��1ネ�*z�JV���1)��c�t1�K����QC��d=	N 'ל�3�� G��c�O�KH�<�~"=ZB!���y|&��`/�vZ�)$d"�Sy�B7���J�Ѝ�@ѭ��*��`*�9[X:n�i-9Ҝ>��,
��Qi3`I��0�q��\z�&0�t-�q�P�}�W�9ڠ����2�Gl9Њ�Ɨ%b|��������� $�V���-�g~��"-��Ax���D��S��ͮ$4~`�IЊ����a�u47P���P�)q�'�˖1c�}�?�/ѿ���/N_ͧl�vF���׾2��ˮ%#��Ӱ�]
T%�H�i�/!��[E����#���l8�,��?�{�j%v��c
���h��{�~~H��'�������|Kf��:�H���RBndIwя	������0LA+�����$�
�����1�b⋉�'� %+�
������&/	��9{S�s-l�!K���5'