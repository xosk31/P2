XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��=��ȝ�ky]�uq�}U0wT�?�5�*˵�dY���2�N*�)J��J�(��7���'~��w�30��}���]m�!
��2�h�����-�;x��5��>}�I���/i��pH=Ѻ��i���ƀ�HR�����YrB%��dY�㕷m5��
�+�At�L)+$D|8e�m.��:�A}�|��gAs�*����{��~#�m8#���3"�O���T�lX��^�����-\� ;�?��`㲴X_�	��4���uO A�D9!d|1U�S6�3Iw��8��['r~�ֆ�*���W���~[jļk���k�7��=��+9p�jG���	� "�-��|p�]3=9�������
�ǅ�NHA��}i|\ �|;��ތp��Ԩ^KsA6t�)T���a�xwӼ�����8�s��U��U�Rf��3��x��9����",��V�T	"1�ZiTE���L���6]���8�⦚B����Ħwz�SM��0�o��S�HI�y{[�^��5����^e �zc�t�[~ϸ�&x�pB�Wtb䆺��OM�9D�}��a��o�ma��R�*���&cU��Oؙ=m�j���}�-��?�1�Z�#��C�9[�y�{!O���.p���:A��9��6Y�B�� ��2��u�p?�j��b�^̮����mu�{X۫�E�ya�^��ݻ%j�Fol%�%�!�a��[9W!���9q�/�j�J{�gTd�$	9HHa�XlxVHYEB    fa00    1790���U�F̎�J+�D��l�������WV�k��V�TQ�ܝ�Oi��fc<�Mh�]tɺ��V��_u{@}?>
����t#T�1�R�z�ί:�ot�Ϥ��s��k�!\?F�M��3�-T�`����Wzq��;��6�R�c�BE�|�pn����;��t��t��w
v����SS�^P0g*��h�_�l(5nyq|������yi�������DlDĚ�zQ��[6���m�M�_ q�~k�q$<F��I櫹;�s ]�V�8Z��A�ZB#rN��.�٣
Ҙ���������f]6�Q!Td��~]�7�LsvK��)�+N��fv��3��?r8�zUvJuɍ9�t�>�Y��`Ax�r��4PL2l��~)��ʣL���&�F5�.,�Ŭ{Ր��&7�,Wq�+����@�mK�GK�9��S]�d5�5|�S�]->���v�M"F�b�uLW���I$���
��WH��vcz�xP��uO��A��OJ��?N��-8FNw���$�����h�͖oź�,ރm��'��Kh�+ �I�c)Q��SI_tP�V��
����.c���34�»=I)n��^�p��b�ٞKLZ��ى��!�-�iT��9��o���sƨ�� �*N��97���6;L��,ڋ'�<�'3>�Bp1�}	r\/�2b*] �Ӻx��'Ä�K�^'��9��.[/"�'
8y�jfH��*1��N��I�J�Z��\�����K��}wxUg��bp�˫)�]�M��dd�*��1ea�#�c�������VKT�n�!���v=%�C�#���6L�ST���c5'0%���a끬|��$1�e�tw�8N@��IO�c2r$�N�j�iKl@�P�DXk�3*2Y,oh���H��%������}l��S�{� �9�vk�fE�'�]}��HԪ����m0����P0�'�s$d�u��Tz&rG+��L�m1���� 5� ��Z�	ө:o��A�2�z���!$��B���X���g?�sO6@M���y�\p�>MF��`d���a�\��L��L��ۃ;N DH�s�Gj��h�{:t�g�@Bx���)�e��|�حx�7���y�O�gr������ʎ����cw_H���X�ʫKM ��� �_h��d����T�_�Fשh%���.�zg�k��D���O�B`Ѝ5���� ��0@��>�~^!��L*��{ z}W�Zp��)FM���=�w$����qe'˃�љl�����Q�:UCv>�T�#Y*r�g�)Ri�|6�H?���ᡂ�`�s�_���a���O��?dAk���k�3�v�/�Kh��!��/h
QE�^����ڃU���|_I֮fi�3�@�� �������l%�b�e{e��z.o%V�<��H_V�6�c��e^l�;dZYn0u�"Cm9=�v���S��?V���'�7� zͤ�o�����oĎcq^�p�p�B�̜/j+rIޏ<�D��B��=����┠׺�ݻ$��6��M����C��Sj�������'D�,��@|�ؽ2��}bf�Q�������!�2൴:I�w�ڨ�0.���4 ǡ�twx]�U����b�bq��Ip
�9tJ��?t��9Q�rKo&�.����r�K��W�n2����9%�p����r��@�e��Ѯ�m�m~1Bv�~��y���K��U��Ӓ%���}�d��X�`0��I*I-�CB��)vpj���uw褯��.��{�ʏ�=������$�,�d��7�@�}T�B��J�n���\��;���X�/��[|єz*D0Ƹ5ʝ��&O�
�`8^øo���� �1v[�{��������W't�`��9|7h�H	Ia"GJ�����-[��-�1'�jt��O��a�?_�8YG��c'��?�ŐS���e� �'��to��t�_ׅ,A�gD���9	$�&�2��\��-��4w��i�����9��s&�L
�1�^��9�Ԭ���d��Vgz�������V ��O��_�"�v�-��Yc$��	Qr C�p�m�d�������	yuW���GBFdr����2�"��5}o����R�*8�o��"����H�����P �D�����-��ݥ�f���|@4�5��&����á�1$���7�A�x�e��k�$�oa��D.��F&V���� �UYMu���+��ý�L�{�e'd��\8Y�
�j��js���U�	��K�d��"�h�ٖ��ch�C��U�k�3�O'��2"Ԥ�)��y��yUNc>��9Ŀ�����r���AX,�E��HY���ݽ�k!:���邇��A6�!���^��3q˺�K1�2c%���i�y���icw����\G�<��7l�R�|�Ae�T����ob�	yi��_���n
+pϙI��?8\ک��i��Hdy`{9W���+S��r��ĉ��fs�w5�k|Rɓ枿	V�>��,r2��?B�p�BF���[�UJ�[pV% ����Y4Wu�x�Խc���B>�X�k��BѲeX��^r�Nة�km�Ռ�Al!/}�=��n��׼���?J.��H��>(�)���Y�W�OB�v�jii�(s�I�� ]���H�2��0d�x�:�Wq�11�r�*d����>���A�vz���q+t��%���yv`
�2C�a��#d�i��[Z�-'.`˫M� 8�m�Y�M��u��b��`�4����`KCgiE6��͕�Ur�RL��щ��+U���+��;�{���돳ax���`�����b�\��TP�Xѵ9�X}c��a�
":#1�UA�{���ͥ�ϧ���Q��L��|�/����D�y�z�N,r֙�Β.`�y1O��8o<%[���;�c�1�CJj-E�ewR��.��^l�/������2�nu��.v�C-,��#Zeq�Q��R�H
�w�#N2(��wQ�R�ɀ0*-P�2/�Gf<���24v4�K&c����W	E�Z@݀��>S,3�N-�PW|R���U�R�Q��;��rR�5��+ĝi�� ����Ak�^�������0�|'�DR�ɽ�p[����<`pC��M�E�����w���5�-
�⌕_���у7�c�v����&d�V2��*y��sB6�R���A�æS��c �~gD�#B�®���ݍ�;<���2�J�ëS�Nh���'�6�Ҡ�F�8R/
�r�mR"q�^
��sT8;�2��Ѱ�\���q<�8�,��Q�I	�G/�.��,�b�5��9�3_g�_o�����Fq~�[�}���T�ᆿ�yd_���*�s����{� 4e*�; 5��l@��bd#^6�p+`���e(�`����΁����Z'$��Gb��\s�u���ʛO��fu�%x�(����C�ԝY+TS��_��U�qϕ���1��;�4_?�4}���O�d��t� Z☮܌�v����7N��5:��e{�����p�{��P����o*�!���x �L!�ba��ڀ�9���1ڹ�)[!����ITG<�y1�J#_�K�.�W0_�"M��&0�qB���&TR5�e:�ЫfP�+k��� gf.�)Lg�E/��R��0����.,KCS���췳)>�OoaO���T�Fq�����T����3����&��pHޏh�:�i���Ds4%V^���Q8e��U���L�q��q��^���ߨu��cR$�l�k�I2r	�T��a�a��p��!���~���0�����>�W�O�eф$��-˵C̊	�c,+Y�`�!�~'n�	T���o��BMX�页t@�,̅:�F7�9&��,զ�67\\��>�DSc�8����CQf�x�U�A�K1�Ō�Y�T	=����X��ԓPXi�Ap���@���*s�/�T���Jqo�^$0�\����'�?��np�yLVQu,$�g�
�^!e���&�5NY�(c!�Z��>��7��c��F.F�;�Hky���> ��[Os���+auY��<���3~�v������S����h�bH�K�&�-�7G�� ����������N+M'���9[�g�9 ��i�
�p�u͍����9��� ���<�T�$t��XG��Bw[�\=Ny�'�{�1�b�x~
��C�����\ԟz����&�LR�*K�v�0Y�F�0��b;TaR����{����=A<��"����n�M���4��@$���k�+���Q)�:�<2�o��yPɀ��
�'"��D�^�=�U�GВ�tT�gM��+3$�z���-Gxd��B%���A;p�䌮O}��vRr�q]���$8�H�jݥ�TLF�f��*
�=�OWֶ��5E����k�#�c��P��R"h���=~��J]�-8��?�FU�H"���O���9�8����2�᫧G�j�Z���.�(�}�5��5����1����_���?pO7Oڐ�O5�LqZƫ��I��^I�i�x�wo����JUHf3�`÷�Ʈ�x[�~��@���^�5���&'�4}R���{d�su�����3���]c;c�]8�(�؀��=#]3H�3�g��ψ�DJ��c�Mep��$����׉T1{����6���q�JJ��R(%�Q-�}��y��)C����Nf�m�H����u�'=������<�����]�ه��lJ��"}��݉&ȸ�l�2NTW��P�(�~ϒ�Ƙ�)�<y�٪l� �"E����A�q�@�圂jƕ�T�D��qA86X�'P6cO�<gcC�I��D�ɑs��X��ʉ2�C�U�cIu�tYy�V��h��N�\�o_df|۸>��B���m
%�E�����*�&!����6� \P���d3�ǌ�4)�����Mf��on�=��፲Sx"���{��nA8����P/�~�6>c=��c<�զ�K����ŔT�������'���Q��lX�{Q"7�\E��Ȅ�	௮Uݿ6I���V&�z���W���ۉiT�jEI���I�U��&��AC����в�=ZH��3
���$��)*��kbq�I#ͦ���|���l}v\��J��,��ic8���$Ҡ3W����ɳ� ����O��������� <�i��?W��2�A�9�x���j�gJ6.�р�D;y�*齤����i�׳{����5A�>��2������N���"sGNR�|Ǘ����[�����jV�09�q��dPd��$�L�u�5{���}b7K��������1�8��X�$T��-Ƹ�u�::jɀ�RvY�J>X˸����MCH����Pc�X!u�=3�w�Ȍ����q���P*#����p4:��6���k+�
8�b��1���뿧���-�N'/�k���5(�FO9�k(�� f�Qt=�zf�择��*�.  E�3������W	�N�[��#gi"y!�1&�۔������hM�s;`T�sr�ИS��������'���SǷ���ǒ��;A�5YJ�7c=���l��cy�5tg�Z��i�iEJ���|�GX#Ǖӟ#�A��{
�Mȝ�>�rQ��4�N�I���e䵫��d�Y��<R�{�L^W��J�	qI�ζ�\=Pᶙ`X>���U��Vttn�����4�l��4��e�O�T����'Q�"!a�1��D�&/���!l̈́]B7hhҤ�=��gML����O��0���5�H�/u��̈4rCF"C��G��Щ��7Üh^�Q��1_�[�S��*r�^�Ĥ��܁�l��%�����~(� ��A��e�[��f���V
��7�CE��Ȉ��N�"�R}��l�;?�ku�&����s�����}��~:K8\�%�r%9�8��(���S�)�ՙ��XlxVHYEB    fa00     5d0[6����7 �-�i���q̗�������0� '7�bˍ���O��.m0 ��� W\���7�����`mF0F��R��fl�B��]��M�����\�3�GKg��Nq���ߘMe'��E�_�r��0ZQ��}Ӯ���e|W�{���ԅ���=P�Je�kS'�M;4����#8��VY����'���Y�i��'�-k��?G���ɭ����f�ۍ�"}�=���1S����@J0�HZ)���1f�Wʱ��z�P��
���y�����W�e;o���)3*����^�����5��y�V��
J�(��|���iO�A9��ǃB&[��F�#2�T�&Y��Fo�@o��-Kz��A��Ɋ�-��10�����+"�bp���)1�=w��@'�ou܅�*�E&��	ۮ�*��U��f�U:~mz��)R����T��/���Z>�j��ӻ�,�l�/Ws�	��W|�#������b�93 (R�f�4uS�~��t�+��@��14����I�pz�9���g:b��z�e�P�uf�9F5W%�ٕE�/q$0��f��R�<�`,�~K>���������?�h/�۬2����>��	�D���=� p�jOX�J��\@N��I�%s�$	����~Ƃ�GWn���?���9s<	8�a�`�G�,��j��%W�������� �ÿ ��:]w4իw��n>m�q��c���?���+�s$s��si��̏Y�V�O�dke5N̈́䎡Mv?�U�&��d'/�� �x`n�%�����*ܺ�J�3} �O���Ϗ�p�4Jɧ<֯:G�Z�,�2B��������{l�\�vˬ^�����x�D�'v����i��|�_mu�d�r7� �F�/�������(�&�M��`ܚ�y�2���*�P�n�a���r��Xc�0$�da�T؇�3�ɾ�[�ȹ*Q?�ݽ�d�#�C`�4G�D�TLu}{����6�cb4,�ǆ��ky�Hx��֌�����<R��k�&&:]��%�r�H�9a��TV/�-q K�SЦ��8ط���X�1�,�K�wd�̈́#ۮ�*�q�ce�M\l�� 	��V�
ͱ��Y/���vXz�A�~��G����!r�¬nz�Q?e�'/}��^y�����X+M��J��"����=@���0�2��ş)[K�]��<���)�2#K����J�_�1R^|�Nkn�ȑ��"��m��ߛz�A7'��/��䜕�Z�ʐe.��>� ���\�2��2��_�����|?H\���N���<���u�2�Ǥ7���?$b�)V���J��֠�̛o#�l�Y5���O*���%�h��|�`�V�#�J��iΔ�Y���sZ�L%5��a��hhrCqھ��!/�T�ICΤ%R��a7)z���P�Dv�ա���y�K���N����g�(�����$Ʌ������dXlxVHYEB    fa00     640Y x{m�����(�=��Zhk\��5j�������S�/���M��Tџ�2�Y�����ڛ�!|I�nL���W�Sa�n[�x:9a���c{�W��N�Cx<��Y�è(Q�U���yJhc����2��q��v��d7�dN2f!.��8�ԙ�� h�ݽ��>�O�\)���`m�j�De�M�dg�X#C���$@Q��CM,�@���ic�� &�«��iBmF� ���r(�ڂ���A/���M�'�yN��ڒ4Ca\����m�i�$��7h}��I.m�~���2"��.�m�����C
�~�	���tQ��K�=��������7>�+z3�l�l`4 ��h���}q|\U���0�}4�[?���(��o����Ț���R" GXv��cc⧻r�T���K<�8�(�ն��!z�����U��F7A/�^�[R���+5�ۂ	�L�(=���Ȫj�-!���}��<���)���0�l�Wv"��W��k�f��"�]	̡���,����k)V(ٝ��8`Cjx��I�a08�Uu�� ���_A�|
p�w{<pޝ-��+J�&����xC���;Ŷ$	p�CLIJY��0`>XȌ� �1�mK��cƳ<���Vl#fi�Ǆ�=Z"ݯULW���@�_��F�S%�*�*�)e��[ق^��kN���p.�o�2�K�L�)��� P#�d���]����3����6j�e$ �o�=\T�IG�	1�6�^��39AV�!П�������!�d#A-�@tO�=��ڮ�jm��Q3p�􁤃ٿt��$�p���؀�L���/;3����N6��5u��\����iq>�C�NƟ������ͷ�zM;}��	���a���T�F;���k�穼���������ĉ�\���QD~�?aMZ$������;Q�|I4۪nPΪ��w�
C����5�����6V��������1�Ovga�\5�t8�Ab/�-�/ɱ���	�0���v�5��um���|�.]��P��Yp��ׁ��$�ؠ���4�g�I����v$�
N9���͡�5�<�ED�e�˗��/�X��t��<��	6���,d�Q<
{�f�s�&��@��/p�s:�X0��q`�!߷�8۷�ϟěO���Ꞙ�R�c����S��l��\�n�K�o��3��gawL����]v�����&�0��3@~�Em��B�a���;%U5-�<G}v��Sz2+�9Cq�l,�f����	{�gb"�L`
��ĈHCS��!���0`<�Zg���!|�*G�
�X	�'��f��O�|�AhB*c��ȼ(>���Wz�L�p��(6��;�I֩G����^#g;oe��l��@�""G��4��k�y����6Ȥ��+���\&|ߍ�R��햙�0���9���t&�Յ�%"���ҙ������>�Y+}�� mo`#����K$ˣ�'F�h���������-���P�����h&�ժ���%v��t� έ�rFA�uN�a�D��zHzP��#-���c�����'i�XlxVHYEB    fa00     5c0���D��	廍G�����vcwh�q��� A�����h=��C�bS�M]P	�4�y��<K-�f�\�p�\,�V(iBUW>u��c036�Սk��w"d����q��l�.��k��цKY��ohN��Ҷ,�������R�$�4ˮj�.���(I��ڞ��sG�}k�'�^vh������-�n¹���h��޺\�9��#MyE'�3_6T����[�IK$HV�T�}�W�:��.<k�<TuPT�^4R
�M�񎌇����k*���z�b����Zeӏ�0�	"XW�����k�$�j�%w�L�w^�Vda�qAy�7�=�e��N#���a	�;��n����^�������!�7:p�� �"	���?�tZ��@ �Hνo%ՀA2JC
>c�S�a�-d��oD�#V$�ԛ� �y&W��3�V�>�rA�{��_LT�V�2c��п;���4��J
�;�4��=�R�pG3��	��n�y
\�K,���u�2�e�F��mLL|���a��u���f����P��b{�D[�|��i�z�@���y��E��=0�qp��*�Tp��<X2��zh��݈�0��^n螯6��8�vz閶��.Ȇ� �,�5���~:=C7��C�ڬ�`zm�aG�ķ��
����d��N�6�Eug��v���U_M�?'���@�!��d '� ��[D$q��^��Uk�5&���i�Q�pF�i5jc�Աc�%ݺP|����0���hLu��=�+�M��C˕$q#n�3?�V�V"����|L�,Я�10���� ��3���c���h�'�'�0.��n�pvTM�`�(�W���?J����ȩ��	ޯ ,��d���ߥΰ?t����L����^� ���ʏ��W?Gѣ������=�,�ma�G�q�;K�
�j��j3u�
� $���5�b?��ţ�{"ɻ�4�Y�=�qa
 D!�=�&��+X*�FcBr��HA�kI�<���.���;�Bb��<@2���?P*��g�����o��V���$#+kU�� �� %5̀2Y�[N����?�S� �PSC֍�쑝����~ �P�����P�DgJ/���
�����d�|����	+���4��i5l��������<кu�������p�]��aRc��w��?.m��4�8 �ڸ����#[I��e
��⺗0 *k�����]3#4�V����Zf�;v���i����^g<4� ���f�� 9��.!���O=޲Z���?�l��%o[��Z)!��k�tԎ.�E3���~�'Q�o	�p�k.ji�탡��Rn_[�k��@�;*j$�+��>�|0�~0X���e+�:�4�WA�U�w����D^��&tL�)U��Xԓ�QW�3kl��J��3s���.J���3�w�B���x̉>dF'�XlxVHYEB    d347     a90>̚H��>�������Z�t�����v.r���9|�cI/^��Ʋ��	�P
�,���f�a5{�l?/F7h䟅a���°��M��&b�������W�`���ߢ���s\�@�s��K&CX`�:Gr�4,�釷R5�v��D��~��E���l��0��t�KP��]{������};��B���3��*��q��b�ِٖ�l(�smI�9��,��J�(��� ݳ�+��>��.h�w[�`�hLJF>2
w���dӗ���O������p���@�hƠ��foB�NZ��%t��G��B�b����{��͍�X��}.1~8���4_��I(:O.en�}&��,�����γi
��7P2g��K���o#\��y�ɉ4��w�>Y'�&(����ﻕ=�A?Z?�X����7̚��`�b�0���c_@�/&��LGݮ�'-M��8�`H����:|���[�ߵ5�e�
&*����QVE�xg���w�Z,���O�(�s55�蚜|��	b-T�|дPS�����V�8�s~����#` �����ȵ�.��F1��jZۥk�v��0�����'k?�Nj:�@�1B�����n�
]a��i"��"�9q_�����4�Ρ�'֚��4㳜+7����W�*q�&O<���΀�w�1I]��E�$�a�����0o���f�R;��Lo��?�s�� g���}#c�>λ�v.���{g˨Tq�&����췏���R�kI<�w:�/�u�b�m�D����|� _ �5T}�ǔ1��d����mLIbɟN���)� ��_��_xBx��\~���3��O���[ͳ}��;�~_)E�8~�4��ٞ���%j�P�d3h���1A����܍j��ݲ���beV1ny�a�0)�ۛ�0$k������+���o�tA��`�c�a;�-���84�lӿG%�:�I��i+cY�{�r��f��ő.j����kQ��b�d��i�lLz~��kf�+6��21׻���������)���tv��i��}�l��t�/	C��R'O��0��� �\�\�y���A3�'��R���݋�8�$��31���F>7��kz�2��)����u+r�+=�� 4��k 16ga��D�%ܑG��3Ƃi��f���2�L�ZQ�(m��X�1�TBq�n�ڇ��6U��ު4VA�Ӝ�.��"������4�S�-l�8�%��� G4ʀ���u�Y�aﶯ?��,iX��gY�%k_��iGV�q�|�e�oE�lpl�`O��Z�ߒy�(΂�Y�+;!6�Xգ�>��ئW�;5�N��[d���H�y�E��֯Uhk�wVdu���L<�2��
ڔ�`��(S��T�s��U�-��E��eD�Y��b@�I����{:F�4U�rA|�q��jCn��k�����=���2~"S�κ����*��K>��֮/�Dȇ��_��Qc���"�_�WAnj�9����F�~�@��d�v���6hPv��M�H����x��$�0��1&�\`����,Yƚ��Ha��i����cb�1�ٯ�CmD>���K�:�Xw�'FP�}�~�ND�e5���)���2�{%�ѮD>��<�g�/a=s.���0�K�<�ln�熼I����6�\�d˟�fab1���s!'��ߘ�b)È�!��Z�p����K/S��I���$��ـ�K��n�U�Dq��dੁ۲s�Y/�5��o��sI�뀚�'�OGa=8�E�0g��1s�|k�s�h�*V��n:%�[n�����^���Ӿz̕�bU������X��!��e��ʻ�|�v8����ȸցZXnV/�+.�YBm���Y���Ӊ�'��h���x�l��u,�?��rT	>'��G�SC�v�~]��e�]��N\��q�:�'z�yު�4HB��# Yy{�b��L��I�|��P�?2���oym���]����JVx?�A����ɕ{��q5��6�'�~��y��U���/����y2Z�ń�u/6�BXo��PmE��\���̋�N{\�r�\Y�Dk�n=�k<шA�E#O4�9��K� �PƄ��hF��|3㕘3��;��;L&2���Y��"?Ɵ��Q&d�I �R41�!]B�ٛ�"��wx<�[só�&1Q�0��6�M��Tp��O��H��	�7У�Dg�����#�<�@�ч��q��N��%�R���F�nl��H��8�����"��_|�,���ѿP��rJ }�C&�TaN9u�Q�f�lHo�������#����� "�E�b�"���֒�Ck���K�2�7�O��`��3�M���֎��mI�����,�3Zuw�&8G
ӆ�����h��p+ �\������b�ǯ�DB�����:��w��!�Z}A7�I˔��\���7SiB��2�(���ޢ�b?���Cc�@��b7V醶vW%B|Ȧ`�|��T �o��v�� �㹞�Շq"E��[E�JbmE9�Z�ol��u��{��L�Q"_��s���?��ݖ|˛'��m�UDTQ�d��w<x7���d8�i8�E�;q0��)�-/Z���=�m��07q<B8����,���6e�YN��x���