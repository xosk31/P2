XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����X�V>����<l*�� Aoe�hv*�|��x��ޚvr���}�Fc 6n��j��N�m�,/�gG����i�#a�������|��{s�D+�!�M�m\ݴ����a���Mzt�^��s�c�XO9n �FF�bˈq��}<Bb>x��s�[�u���\���5�T�u��K��+�z��#�� ���)�,;�U)�u�m*3�ǌV}�k��j�#aI��gا�Q�\��n����*'h�1�$�w`K�F
y'^��(�?�MY/jl�0��g�$W�E@����vS�/;F<�m^t��|�g�[��r�t;��g�/�� �A`q����1��x}�re��>���˽z,��(y�4J#V>0$���n�t���3�5��s�8XA�0���0�����	'�Pmn�x�!z�>M�?J$���r�����$c<�f�R4����r���3q��������]�
���y$��$ ��?��3�����[��SKh�I}S��R!8�v���Y�{(����G��y����L�-X���iԽH��'�w�W��9J������0����E��wXk�<���i&?��)��L����!n��楿^+T��u�{V��d��{*��+Oٟ��[��t� �zq�tZ�ɘ��2��Doa�"x���f�T�q����X^��Fߤ����5o�E�}-�Ǭ��f>�E]��j^{`��^�,Z'J�8N�b�X�l���]͂R���D���diWd��/DP�	�=H�XlxVHYEB    125b     750f��s���)��`�4�<F`'��o4����儐�*�eH]�7L��l�sm�f��͆�jgR�v��]��7������F���X�Wʢ?���2+�PwCB�h5u�T���c�C��k�����S�E�Tl� �ִdj�_��I��u>�=MB|)�6���g�;,X�N�L�
(�/}�\"�b�f��վl���Մ����xg���)�t�����v�܆�!�ư���%F�)范.{2���&`��+.A7cl���\�$�F��h�>OB�p<�dv
&���N��n`� �]ʑ����8;
�fPi����ƿTO�h?��4��{(e��!�[�|{a	���fp�/rw���A�E�1u�;���M��R��^ �g(��zu]��+��Eڲ��q�R$ �$�������_��R3�K�ڨ a/G��n�����.۝�^�FU�C����$��&����O䋔�UT�,��q��R�t���X�V��\�Bk�������(���RcM�F����喎Ū6qLv�?��Z������j�/B���Æٛ����~ld�o(kA���b>N��k{�d�$_~��"�p�hb�m�l:����ݗ��Eǂ<:W��s�X���oJ�Tt����p��V�ȶN��i��:"�Y�ܔ����	=/U����:�OY�#ㅤjh)� M���Q-y�]���`�-���њk�[�W1WX'�#���3�SeMMK�������2�GL�cvHu�ϯ�ó汘��Ϯ�ں���$�7ώ�����\�)�.�E��U�$`�-���{ᷓì�<;p��Ks�"� 黕 ~7��ew�����d�}h}�ؘ��P�ԙ-�|�C��*�3(i�&��~Y���<NO��rxF��5UIg�@����2uw8�XJ�%d7�ph��xYr��)he�n�7�9�ElV�\�3��}U�؂F���߫�Ӂ2E^C._^�n!.Æ�8�I�N��x$��$���+�u��)�-p*Ҏ�z�F�Q�ޝ�ʈG�k`o�O;�l�i���&˻�zl������	:��1x�ɣ�4܅��2���(��)���𐷴�yT�H&u�3���1ʮ}��P�^Ƿ;k����Ȏ����l���(Y�,F����A��:���ު�-����D�	�t��_nV�~�UV��f|����� RF��h��O��� �sD�̥���;��r��I�Lʡ�U.�I|ŉ�C�D�Q[����gV/t�ZX�I)
��y.�M{P�;�ql<�����rck�vM�%Š����F����w�*��ܓR�t�g�E��\��Y@_.�;�����3�*F;|�	��8b3:cT����b8[����[I����A�z	!��� �p�nL�uBa�g2z>�^(���Z����]���wU���cS�O�+���[��v�w6�!X`d�,�=����|���cߐ�d�
(#_�(���u��0]�������|~�NDI�E�j6e��
X]��d+žC"U����W7���pcI�u��� 	��B�*߱���b��Y���h�o��>Xm�R�-@h�`��L��G�üM��U���� �g�+(�fI�I�)V���#?��˦�Yě]�.�?�m��rL�D���)�6�$F�"/����?�c�D
�3�֧������M��҆�"߮L<�"�κ�n4�l��UJ�'���!��[?�E3�d�	D�t+z#��A��zU�Uh�J�#���y���$�������Wtvg�l�e>���J�g��=gsvHL��jb���ӫ�_�	������;�����$�