XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������뗢Ί9cAd�Yb\һ�`. 4\&�A�	�v����Y�v��M<:Z	-!��Vfݚ&�e����qr��UB/��QM¶��c�������Zc���J�'`Q��9�s+$�lɢ��J�p�|)�R솘7�@�����:�"�\�ك���s��c��K�@��.J�B��U�;�K���3P/��g�j�"[*YSQC���E�+u�,���n6Mڪ4Wf˙�9UE;���v> c�s�c ����ӊ6�*���,2�
:������[��!E�f��O�tl�������ŀ��PR�A���( }H�f���&}�e��}0��c��� ��q֬B�T-�Xj�M�7�'��q>��K@u,j"��&:htH5�L'�GC��'��p�����,[2DJ��<��A'!�6�/��OӻB���Fwmf��ȹ/��:�^����%r��Sн۪���;��t���<��t���MZ	C{��P.@f�`��e��#�HT�#�7|L�.�?�Y%��߻���O���J{����i�NR6�6)!���nm�'%�5k$�i����ò��9���E�jxɃ�X�}#�a��.�*���jC��#����Fܿ�:�oF��h����Oَ*����s�H �����w"v�X�}�b;e���&�8n)��A���V���n�D��/�g�H��ܹl���>��v�a�>F�̹�����[�>������p�Ͼ/�T=#����{�u�د�XlxVHYEB    2577     a70�٘Nst<���)�%|U����
�!���e�k�a%�gH*�L�nƔi�$�I�Q�c�Q�nD�_�\��;Y���<���є�T���HY����RM(��E�co�;e˰.�4}��-�3ٵ�� ��+	��J:�*7��O�2�ouX�0Z�i[���N*?t�k��/��"��>C��Ƅ�Z(�=F�۾C�GOصr�U{�S;ԝ�[���39k���W\�֛�A,ا6��S��5����g��@�c�}���|��Ãza���(5Q��gi���~l4C�Բ�|�z6&�r*�'gV��5�Z* ��R	_�.�9���9C��J�k�f�������QM�
��ע.��B�i�
	��Wv�q�[�ϣ���N�"���`=3' ��ཱྀ�`�q[ke6y�vH��7�d�BgM�R�OF ��~���li[���!��C��q���&tKSK�N3^�X�d֐~��=>�h_���>��}t*�z�;�ME��|;��aN��@��+�0m����q����U8����u��ڝ�)`���3X2Kdc��>U���~�����; BF��������Q�/�/�Ԍ(e���%i�F�!�y��7.�`? Ψol�3��SGT��E��:�
+K�L��Q"�Dt����|��*�QO��.tX@;��<���:>jZ���X��v�w]���@m�-qp��ʮ���?^-�����5����[�{͇�����R�^yP�)�s2�<��DO�0�v�%s9�w����$D�h%�=j�\���a���R�϶���'j�6�mW��X?�����_�#��~�e�7徊䂧h��L�+��o��#>�$��48.ZK�O�uImӵ��ZfV_���Ln*��S�f��޷�ͥ4>�ߑv�q�F�SѤ&��)_-�!������@��L��A�`Rf_C���#I	�Q䄃�`�]������M1�_��o@n���ٞ���$)gd���0i�6G�S��̀�a���O�#.���ș��2w<8sG /��N��+?}З�-��l���ַ5�y7%��3�^�R�֜�G�2_&$	�͏��4��4��2Z�~T,�k���Ѥ5
��j7�~�٩��2"�\[��	��r����ਐ�%�Aܳ $��Ho��y�&g)�j�,S $1��K��!h�U��ɣ�P��\a\m,ʭzBq�Gp���3:��u�,��^�tG��xi;�����쵣^�_����w%����c��$NM�#��P��{�U���F�� Fa�]�,���&x�f3ĉ~+��Lr8�b��W������~Va<y1�j|�DC0�ڊ�G,���-~�	T8���ALi�`<>��j�
J�Q��H�������_�K�X�P�b�+f6x^��l�7T"���4YJ�X�tg5Ӈ�h�*��d�����4��9,d���B�ͻ���*7!�V��iW���P[
ݣR8;�w�xs��K�⯉�(\3�F�	���B����0���A�L��S� խ��n���hps��esh�|��Ȁ�H����A�E�h.�̸$jlR�@�5d�L����ٷ�]�0�
@��]��v�����	���.^�ׯ���)�Z��L�� bd�����:��9v��0SV|`9L����49�{4��M�	�x� 
��q;��v���6�G �R�F�	����O4�x]�b���p��_��v	IJ]YM���vz���7��,'�Cx�А{�J��c^P±Nf��GW�"T�J��]�L�N��s�ԧ�'���(K�� ��̃Boa�����}azp��cx��;,�L�!�'AC8Z�&�c��xI��R
x���{hC����y��JxB�>�:}���x��{ذ|$�1�O|��tpNKe�`,����UK,�I�A�]�K��6�����f~lj����y��vI�X��R4�#�������Z�]���w̓^ф�W���R��ƾ������`	m������2t�M�5�� ��6��cK��<��P����n���s}�kM)%F&�E��J�E��΁E�Fl*Eͽ��0�Q%��E-��yI� �#KnI�GXMq`;�h�ƍ��� ^N�c|���X��L�)ѡ-�B_??�):�(�-"o~�l���Pf��1�!�Jh	��-�����vRG��=絊f�@���Ĕ�d�c�S�q���;@y�6�CR�"xz,���v�0�t o�Q��!dzr��2t��E������ͻj�1�A��E+:��K��G�i�JU��ɳU�a��bz}���ɰ1&���p�BH'1�'~��e�T[ي�Rq,0ۺ���]�x��t'�2-o�)�>�� ��:�z��\�����}_y��V(c�s�n}�R��Рdei��h,��k.�ۃ�����C�}@׎<�/!ʵ��wǎ���}�:D�D��D^}�2 ���w�ퟶ���h^��V�d[���HUA-���3>��ա���y0w���f�,=
<�&V��O)�Dw�\a#���O�6;r�,���ɬ.���/��k�pq�-���-2��ע����.;��D�f�QM��?�|T�YPF�Hp��