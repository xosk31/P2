XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������ ��o�y[.����)�c�^#��(}i`�ua�
�S��S$�e��:>�O3���b�
Al��O\��U7�
]6��ؑ��W��d(�IhL�f�M�C�ah�D-��I��j54�]����V� =����
�'2Q6\�>��Ci�	�O�9��,�j�BtV��.��=�_�(C�l���kW7?3�l��8�Tv��=��J�8;��g�����N:�;BG"�ǥī�6�����<��-��c��f<�ɭ;^��`f��✕���=�י�h�V�y>��>Hu>��������p]�j������Rr:� ���n�UL��}!��D�l��@ �y�>��Pޅ`9a�aD�	g:`_>��2ޖ%4�FX0�ܥ�ۋ���n(�0�S�pv)a���i�l!n�fv{�q�3��Ȕd%��2^6����x18������W�@z�H��ɲ [��!�%�.$5���G�5�����m"���#��+��.��dU��\(l��Ks��mot��+]�Y$�з���^Y��Z2'�i@��48#;�����M�b��w`�71��d�� SG
�U��'��[)��b2[CwB�&�î<������7��d�����v;� &`E�Ŀ ���n���-i6�Ϯ�oofF���=6Bk��"v���y���Z��aw��������:��yϷ��+�=$��}�-�A�9t*�_�j�Asj#7Ħ�T�Cc�����1cZCƑ��J9��XlxVHYEB    9193    1ed0b���;S?�RF6}�
JڊW�6ws_D��$���8���h�����#)��JyY�� �2����rM��$2R�"%Ʉ3@�o����KPߥ"�U0A�~<�8�o/����y}m7U��P��t��P]�M�d��-��]��&�j@ZS�@�U6��1����L�h��� �#��/��_���Y$\�
P#ȶ�8���~�2z$�*��L����s�]q�{��?읛�z�Ч�d[�9��H��0��Y�m��6�n�T�(m����W�\�m�a�����9V��T�4u����F߼�dIg
מ/"�Ps�����Ғ`Bt�]�g� *6�C�J$J�4P�E;p��<[�7����L"��)�Rvj�C|ڣ8}IjΩD�c))�	s&���D|xO6�*�$��D�!�{I�]�B��#�\yϫX��$�(���H�Aay���M�e�� +Ђp�>'ɶk4���F-����J2��6����3ZI���C����{�D����Q7���j�ɋÒ���M�5� J���
muiǞ|�&6� Z���|#���Y�����VW�k��Q��L��50�%q�V�S7SY��B�r�l�yc�t����������c���)��Y����Hg2�Xe�Z��6B=^����j�����٣o�GR�ý��޸�b:�Hw��Sm%��d�L���`T�#k����3�k�0����3H����5XH5�V=0��fE�*�^ױ�y%)�w�r�˵kP!�2�������r�O����E��O�S;�����,&��壗���7�0�d���!U�4_ϥԿ�\�.T*T�,�Řխ��y}ok,
���E6���N�;��kDx^Ř�,S�ʡ���vs��'�0P��� ꃭVyڞ
`�*�|{{;�@�xż����7��!w��Z��zM�����8�}�#x`f���AL���Ơ\\:�+ }��:�Vphe�-�>~n��� ȱD��e�u�c\�T���c�YƔ\Kh��8݇���۶��Ѷ4<(�Ni⢁QP�}��]S���pKl7�r=��.R�y��ؼ�=#=Qa�_=�no�O2��5~X�_��ڛCV���m&�����W��~ S3�j��$�ܝY)�Sz�K�Dh�P�0��J�p,��]���J͵��%�K��ox�O3;��mD5�	]��A���Þ��揶�&{f�j����5�U� ��tW�xy��C�ǣ6l茤��2xyn��)����\�ix��o6#��%�@��Yg@��m�=�<*6:{]�HPg�� �Xw��h�b9�����]V��0�%]�j�~�)�3���gR�^[��l?7R��<KL� !����#���-�k�� �H;u���p��ݕ%
L�390h��J�5gpјK'�ҍH��t�uѧ�����y���쑥�X�H�N���>����{��ʋ�)���M�4�{xI��l�2ȯ_��>�Y��';5�w�}�.�/�A�9d���BX�.����{�vv����8���!��#���2�6sPW���F�2�iû�1Z��Ŵ��(edz�xQ[D�a�Hsx��F�ǚ<[[�O��[������2�P�n\�"4��>�g�%�1��Oqa -�GbFr�g�p�	1��<z���<n3>�܊K�P/;-�F2Jf����8".4�^�}H��V����l����_T��,0@ê���R���9�Y��"O��"G��;�K7�j�he
��L�p���8��3:~ �;�Zಱ���/:�U�#fr����H��q)��� ��{�W��g�!W�>I���������T��'#��b�����|Ũ����s1GU�01 �J����>�vj$�4�����䛍�R|��
�-���h/oX�d�ٯ���M�T9��a��CVV�$WJ����i��BI��W�R=9�u���,7=>���X�i�=�%ٽ���{ܚ+"0�3Ϗ�W���
 ���o��FӐ����Ѳ��y�^+a�����]ẒYƟ�ߣ.����� �����Q~7٧?a��l��:�q�5c�-bN���.����I>ۯ���M�^F�k,��N}����@���XL��k��KR����p�a-����5�7���:[��;����G^�>��ܕ��3����#>�,D�}X1��_G���^vz�A���<qh�h�+�G�o�]Lg#��ݑo�U$�0>��cT��դp^Ј����dx�}C�'IX�.�
���L?D���*�Wbxk|�(��clN�f>)
��uQ�2|�2�}V�1A`~zX&Xz��ݮ�:�l�߰,2�ך�V!+��i�a}[P~��Z ?N2c�(����w��ґ0[H�	萾ӽ�p�I�hIS�1&/�ا���G&߬�X7m2c����v.�X>��ia�$�@-�lU�ā�	A��J�N���N�Cl.l����zu���`"#R^�@�D��7˥B���6���Hu[yq� �z��	_;�Ъ^�� Ԉ�ݦ����p=��N4�Ѡ�Z��ɭ9{��	��Ĕ'�@�<&�$%5	��'v����:�x���Do.�ԡ��i�C4���<�?W�i ̅�Xr&��\[�,s�� �o���m�|��1��v�[{�m�~ �P��i�f�,��fU���l$�a)u��R{H�OU$h�N������	B��5�<F,�]��w+5��;h���O7X+��S�f�����3O\�y8l|3����.���6ǡ�Qܬ@��ӫa����ʟ���YT�]�$�4?mz���嚋�)NI��rG�c��Ty�J@P�;	�d��2��^+=�C��mj��f�C�cI�n���k�	%���ޝM(��k�Lrj p�s ���q0z�-���q�d��:����H?>��K}�\W�ҝ]>��P
� �D��'�Э��V^L����cR��|"*s8qM�N��)�8|}Bf�JM�	�;�4;��I��X���6��]Kn�[xe�1������
�enQMI��j�	v`�}�~��m��`yʝD�i��)E�#��	�����x�!O��v�Eס#$��jT+y(��|��ۈ�ހ���.��o�c����ڝ´�>��E�����=�rp�$��ʏ�w�$��|��>�1|��V�[�Uߟ�:������-9Ȑj�=��t�f�nfk�����˦�fnr9Au����60n�����/5��8����m��3�_$�{����{�K�����9�J�\@� 	���� �����.<=@}7�x�8x���R�l�4���*�OY/��$��ΨK���Q����.�:ֱ��7#�v�0!lso��Ip���7����p��-:�G�xS;�7s�&���l�ђ���Ơ�L����j��񡾶R��2�)h/�RIn�8x�q��]v�N$�����n\����� ,k=��(��̶"}h��� m�,f��8㚪l�Z��?����kpI��:�r� �O�Y鱂!.>�P�+yx�T�E�#�1֠��o@��LL�����Ix�p��;u=>pOP��~���RM%�-[1 i�_�� ��>\�Q0�
& O-�Y�.��W���M�818�@i;W�ie���#_ηYw�G@q�J�ᣎL�@�j�L��c�oC;���qnβwD����½;сl����(��C�"uL�
(�!�o�����Շ9�����D�+m~�-04:������1�Iw\�1XV��T┖����@1<�M�|a��`�7H��Qv���q�6� �bVAV��ɷr�yT������'5f�J�t[|�y�?[�x�h{6���mk�C�K��(ڄ�
x������m���k�.���E�����Ƿu����O����a��ka1Dn�^&L�x︫I�ض
=2�T����=����CڤƧ�Ɍs�$@|�8���U̣ga~vm>(
aB��#�ֵ�j�jk2�W�?�N�����[�Ac�=G�ԍ��"��Ԫ�T��9�� ��5��#�/Ki/��;��Nk��T�kh,��R\~m�"�[��m]�f�l�dZ��4�2FK���TIn�ϐYj����#}�Ay����0B\jtG�RY1�UB���+Թ�.��������ɺ3�s��B(*r�	�i������c���V�g�G>��x�`^ܷ*^����/,{0T}T�]�#��:����&yrU�c���Շ��;�8@޼ಌ����C����������9٢�NK����أ�)n�ϣ�S��tV�9r8Wb�eB�~�a���v�����M;��dky����+9��5�h r�ڶ���t7������}�@ڼ�cO<���.��=��K�e��p�f�8>����(IT��io��l�I?j�2ԍ?QP ��X��١��p)y!�?<a7�t�x��oO^	��#^g0������ϚwA��ֈ*��~�lR�]%,l���$��V��&U�@�%]� ����C����̠D6YI����=�	��x�"̆H��\�[�Sw᥯����k�+|���'�V����p��k<�~Fs=���w��W�nu�΋����R����t֘em�:O�����U/�J�hنͽ�Ge�"����u���('����f��/#�ճ��~ŝ�C��������)NV3V������w:�'Ɲ��W�~�C�����4^ҕ�9�G��Ì��\��i&������	c2rO�T|V`A��p��j�*L]�x��@���  �*T:%���r���c+цO7�l��!d�Ʒ�$Px�i8,>��d�kE��8�.��bɩru%���x�� @=!.�?0h���5бʯBN@����=Э3��Z�Id*��K���gL׎P�bA�zY�m)�ߔ&�5�0�0�X�H��Q8�j�"��C�N���Y�H V��&U��t*�śy���R�A۰� �8>�j�j�q��ȫ;���vT�i>����0 Lx7GL����0����e�.����"�o�h�����ť�>���|)�Ȕ.�L�:��gY�x�߮L�NGt�p����C���T��-��M���Z�J����E�'�A�I��bѾ��@t�g�Z/��:�h�w4&�`Vp�T�R����g`d �Ƈ�^[. �M����-��K8�-\����� ��5l�5��Sb$��1��{�K&�%�W;�s�ͯ
��j�Uē����r�}A������u
�&s���߈+�^r���ߣ_=��փ�XEU�J���مc�JBƯ�.mΓ�	���m�*�e����K�?�8�ć��Q�P?�d�5�^��P�B}�J�kFUp1\6/�M	��?�"[�ݝT��l[��|������`f�(V:�d�L2�b�G�7���>&�/��%2~Q�U��W���֩n�_�m�j��^��Tu��N��K��׸�O��e���w�P�2,��1��.�{�:K3i�?��o�GYnB�o
Z_���wU��8x$M�%
���Ճ�h^?�FW�HX��O7	�V�{�]�&�m�^�*ԵG��e�����8���3�9�U4�T����v��w����O�·ِD.S��a� "�{�hȌJ9�#�������s�!^�Z�ٶ�;x�]��ͯJ|���;ِ����W2���7��b�x���&T;`&9i"X;Z`.o�ԭj�H���o�8��K�1�N�M�QM�C,�Dm����"P@܀;�r�^;�-�$�G����˛�!m4�^�����/'�"ώv�|.�B��p[����X� -�Ck\|��u�R�Ā'Q��%1p*�W��K�H�i�EP&������RБ�L��!�ފC�o�Zϱ� �`�C��6W1U�1��9$���Ӓ��π\
q6$���E�F	%h6�s^�0L�!T<P��W��7z�y�gOI`�'�����$�c�rq]&��I�>�|�@%���$xk�K]�̃��X����ᡞ�$8���Է���q\����(��4�±'�+WV%S%�V����� �P�`f~EBI��h�h1��eآ�9tO\���}_pF��?�"��DJ���ms����*l��`�<�%��aP���N��-�:�5x�ْc���f�ZĬnߒ9I���Q���Y}Z7S-×�:ݜ�G�*�ᶸ�H��e#�c�S�<@��Yjh�����~&�d-w3�\R��t��!��\������MĒ�� t-tF9ߔ�TSIe�/�O�jD��փ�`x��ò0QV�[���6���p+���:Us(Й�&�eav�X�*��E}�Y�&��2��j!>�m�:��}�����DL��w��ث��\J���W�xO	h2�eJ��T��v�~�	�����}~��)����୽�C�h������>c�*�fZ-&�s,��ԭv7�A�j%�1k����"'�ܕ������״g�'�vy6r�_������0�	��B��y]EbS�Pp���M����ʱ�X�@�?��_���:�ޟ{��M/B��v��:}�Li[�BD�	�������͈愄�B����ˢ���H���_t;Ȍw��CG��e���.>R��Z<D���O(�	��H6��LR��#�en��홎��P�tE�m
�j��B�b�7�{�,����,�������>��'J���Uv<� �!�wCA������`�/��t�(�`nl�_�`<�r)����#u*�s����C��rE���]��X�L�O(p�{�|���:h��v����u�^l9�=�2�O-���y����p�4�{}��C�������i٢��DS�Ү����[���v��v���� ���n�w_���&���|�������<���v�Y{�ǜ{#�(�;@��{�@��11��ZU�����-��s�ω8`�VM�aM��xg�o%2��m��� D�/d���-�Փ�4.]���V�4�Zh�a0C�}˗!8�X#w6X<�fL����U�e?¯(�S�ډ���oʡ�?�'[����%(t�:����t��=gö���9i#�V�dΧl�b=���u�7�?@c�P��Skm�$(�d��kh�U��E���+�3��p���y�U����F�5�KW�����~Π�L�,��g�5�h���5�GY�&��� ze{;��h�G	.u�H+�ڭ2���ќ�����\G��X�6f1��yA';a ��~�-�`!v.@�� ��\٠qT�X[BL�����w��x>�=P:W"6N���6����_sw/�T���`T���0uG�4�Y�֑W{ZG�����(p�fOR�0	c�jH�G*�I�>\.�!�t�����n$ Gt�[���L���f�-�D����H��؟�HڜS!��g�ջ̫��m����Ci1�>�'��]��� ӛ��P�?�(���*�G��=T�d0r�;��g��%��?k�FM�;�@�y�C��>-���֯mz\n�OY�c[�O��5�e��@�hkn��!{M�y(g5h�{7G��[���:� ���o��_	�3�8�=C��n����|t�ڷ�:N��E���R_7�P�0�AV�	h�Q��|Be���#d�`�w���%7P$�5�"I�λ,��OG���`8'����Ѳ����.�,h�>�V���Wu.Awو�p��	����T�#n�<J��l'��ĝ��� �X���_f���э��