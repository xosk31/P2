XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����w|'}�/��ԨZ�� ,�#�yi�5Aŧe���Q{�g<;��_��B�ẃ_߶7ij��!�;�c����� Jp����$����C0sZK�H����h>��i�k]��/b���xa&C��\㟷�xM����*D��._���ҕF�QA������w���]�&~�u�F
��S�q9"c���OJ8}V�i��&�I.���vW��-4�#�C�Vu�V��q�)Syo�1�>CM�$��ǣ2�{u�"���P�N�t/��ڟ�=��+�EGF�s�΢RGH�SK�� �i�Y+,����+���C�]=�̕ �C!���@np ̻� ��<�F��<s�(��E4r�7YѦ�F�����4^N�GUd�����OK����2�4\>�ϥ�rp;$��R�_95g0e��9k�����Ё���T>�󯹜=�0�+D���
4�tMRX|��ǳ�e jF�	{r�a�2��h��3H�"���4��19�x!٤iQ p�YȒn�)�O�l���O���f�~?,�=y����JlFy6w��v�����)ʾ4����a)X��ǐ(��\�$G��gU����QWj�b��g�=0�����ko3c�G�'WdwnZRoe�g�>���A���@�A�L�h�rG����Y�ҵ"��{FG�ڗ~pA[Zw�|na���:=����>p���w��6qH��6��ndg\���ށ�q.�5��I�4���N�.�:���B���]Y��a%����7�{C�x@��_��XlxVHYEB    4192     dd0��j�,9y^�����E�)�X��n[c!��w��ϳU�rHv����ZVܖP��x����\o]���' '(7Xۆ`�E� �2 H��t��G*fK0$��%�����}�e\c�]'��N�mO��«DqOG��ǰ�̮{!l��k0��Z(���ޒz"ǡ�����@į�����,y����قk�j�@��o�c���G� `���#$%攟fI�V}�:(�aߛ�x��t��r���gY�J�&���[FH\���y$�p��U���t�&�;��(~�;N����w��Ƶ@�����8�	�oU��.�\��1L#�����9$�]��yd�.s�Ҹ"�C7d�f�G�]�s�_���d�q�t��V��������=��K�}��JX���K�j�}yl2�q�,��џ] �'2:��0<X+q$圭��������u��in_�|-��U��wa�b����S�k��=���<%����],�+)�V�e�"A����.����Q�Aޖ�<�S%_�㌝m� �7��Q�:�#�,���L����ι����Z��\����!�'M�S���F|+޴�]�o��!�)�]����Z���d�M�E��p1���ӭ����kz~$s�λ����j�H�L�u��Rm.?XP��g����GP���j�� �g�FV@���7 ���K�yKe�j�u,��@>Jh�w\����-��T<`�{)�8S�.������{`0��?�yy߷+DǢ'D'����:RCQ},��j=ц�X��:)�R��@�K���aX��܅�IL�ܮ��:.m&���)���&B�'`x����Oh�����35��t��
�v�)xm�(��_x���u�oK��.�ռ��7��ƒ�+������w���zg�F��N�x�W��Gсe�|�%�����������ĕJh��"�Yr9�K��1�Nm#p��9dc��q�JPC����4��-��C��i�6ǋ���� ����P��QL�rr���?���t�I�J<���K'9�%���?��Q��_��@b.k�� �D�:�bG�E&�6������YJ�?�����gyc�����^������x�R�H!�+A���h���Q���|�(���H�P�@H�.�'a?
�j{(_���،�}}޷�*�;�KI�'�}|b0�N�k���~B^��TyJ���b%�p"_�q,��=is�����U`�w�mS�,�����l
1*(e:2lM��ڤT�Ȯ�d2��w�B��yhqA�q��M'<�f�p�VL�>E�<����븝�dU�t�x!%|�mEm��WJ�R��nZ��<�9�T���O�.�(OO�0T��B�cT���t��%#��)�����b|��A����\���1挤( {���[jVz'���m��_�$����.��K�#2Rc�̬`�jU_�P1���mW�~���ߨ�7�)�%q-@�cY��d���R^�(�v�����i��b	p�0rWV���@���=n�+3�`&.��f8��4rD5F �L�J�;��9��͂Bϝ�����=�_͟S��bBϱ��I�%׭��2�v)�veO)5:a�@��+,�Qm��zFS�^�)���4���>y���>�AGW�ɢ�T�^ᤝйU6�ϬĽԾ�'n1�͇����p��l�no\�Wt���Qb:�>�-�S'C�tf�e��3{�&��5����P�<��z�0�w�y�wq=�r阪}��qƾs���]�a�`t�j����-ht���)Q��ߊ��Y7$",p��	uhCvO^J��T�Il�چu#��Y*�����"�@�}j����d*�ƘRG���E�@�����'�.�Z����*'2����>�X��G��jV:�%�M)���=���bYECU���"�i^��W!Z���B.�s,S[�9v��
�!��?��[!z���,�Ly���whQ=�ú}̎���F�5�X��?[P��UҸ{��wHս9P���h��;9QU����+��~����%�v�\_����'���R/e
iNX��7���Ma�h���Jp�+�[u�!�5ŀ� �Qv��R/ꭷ�Ow��W�:���o�*�G���ve��G�T#�����C�p����y� ic�>9q�=TIj�hp
�$���wI)��'��$�G�2��D~gD�����]��W��Q+a�X���B�e�.D$�(W1HǛ�����.j���d��deB �6��X�����f�3a{2��vQ
��GD���K��H�f��j<?7免0v���;✔;�S���f|�����T.��OW��ƕq����r	�N+"���Pr����KYb������]$�
��[g*ld\�J��,��Ԑ{D�"+�:YMsJ'<���Nig�P���"m��6����_�y3g6� �\u�V�L.T5����,�{!?I��lu����'��\gq擨�)�}ϳ�l(��"��e�i?!�Z�-�6 Ƅ
ԥ��K���_۳P^��F�[���Rb���щ{�{��ur���z���%��c��0�+</T�e����n�b{		�93��S|k�8�usSG�$c�ї��F��.ӊ�)�H0P���.�����H�}5�i��a�M���N�@�*�y���-�H/��'R����d�%>�iDޗGn\�ܦ?Z�����#�&ŝx�������F��J�29�Y�����l����x2-�3Rv6��k��s��4�2:�W�"���d͌ �w�a����aKr�ˣ�}�����m,hv[���;E:/Ӷ��Ώ�9����������f��/G^�)���[ jU~)�'�j�Z*�ɸ�iAӬ�ݺP�| �&�;����l�I�� �6��~@47��ͶO�U&�=��[��uYF��ȍu�'�O�M��M~�D���z�j�-b�ͼ��;3�tV���j�hP���@�s�?�.&��]b<������:ORV��V�?���v�#�����>�|hq�耆�Ht�X2�p���'�Uأ�ǈS#Y��rw68�|�ʡ�{Md�|y�ۤs����ԣF*ˋ�W�B�o��ft��$M�����Qʹv�q�bs�6�Ҭ�p�_�X��!QT}A�u�� &m'�8j�QV�|.����6hႎ]{��� ��v�MF8lھ2��
�����2q,��9��$�;�,9��f� �J�֞up��f�p�TDd��%t�8Jw̩X�3{w*��ٴZo4f�u��v��Ո�姱\B�T)$ ���a<�R�Om�al}�!Ƀzx#��̞Җ��n)�m��m 4�{@+�hA�{w)�ճ��UM$�픣R�Mfz~\�J(_��0�n�LP^�/�j~K9�c���i;�(�ՈL52jޭ�-����B�9jc{