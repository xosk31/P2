XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����+I��B��{���m�x��"6���!O9�W���Ӿڦ�z�nl�ݩ&ü�:Fm[-� |J=Y�D��`��3���`6�Q�&c=�ӳ_��<�]��H��d|Ukԁ䁑7?B�Z�k(��9]���5�	�g�6ɶ�s���P��%Z�q�iu�T��<�5��3�~���f����L���ϸ��^0&�3�w��\|u[�7Q�%�G�l1{�C^lB�|w�α�U�Mh�D	�+y
=c����W+�GZ���_��j`1�g�����|���w�gT>��a�w��I������\���M�0!���v���i����%�Ґ��2N}س�X�h��Z|[�t���wPM܃�4��/�2Eu������V̀��(9���_~K������7e�*��M<(�H���l�5tE�e��V��uٺ^ќ��tw��a�Dma�Ô���!N���M=\�l�r��u���B��W�{�Y��D��k��U7qM�x�r#�S�6�QN�+T$Yd�<)!���z.��VO��@��z���z/��8FS��2֨�F�j����q)>C��Q��6dA�v�����M���Θ��M��B{f�	L v'7 �@���������R#nU�-B+��5�4����؁J`�e�a��f�PP^5@��5"��&OV���1˫�@{�me�*��<�-�X����,���ES�m�W���Ϛ�`���ż���\�v��@^Z>���u�c)���Z�#XlxVHYEB    fa00    2030�h��Bu�ʃG��&ȼt�t�W���	����������D���ى@��[��ѽ�]\�A"o]� ���0����j�^\g�y��Oc�Fbk�&R�ӷ/Ġ��G�,�2�:�B�Փ.Ԣ�[�6,���ʥX���
`hG�U!eTB7�ᰔ�8���ic����ϟ,��p�R`�P�_�C�W	���ۙ�0�hW��f�<��~N�����8r���RIy�O�\ϓ�=%kU�L�[��B�:u�� ����n%ꖪ����:Z�>��I}뾑�f 4^&��9��%/�VƗ��X@�I��r��xHN�&&^�_��U"���Q�ݜ��u���|"c$�t%:��:56�%��Ę��	�*�m/#�̧��g1H��}\��,�c�F^T������A��!۷����>���L�������N;j�p>���"�(س�l�}����\E5�)�H�>t��Y$*��+���3�?R���1�.!��ep������T���Gm��-w% ��S�#�o�C�}��P����b�aX6��,@D�ũd���"�c&yg 1KU��3�O�Bٵ���v�4ETz"���� �[�S==p�8��{���,�������о֏D{���QI'�Tcu��G6T�!�E��h

1`X�t�M���_���k�e���������?i��5|j���6����~ʘ��P,����5�,><,��&+56 ͅn����>k+�K�S��$cQ����I%��ր��%!�}S�k#���
Ѿ8m$Nm�W�Cܓ�}Gw0J��n��U���C65M õ,��b������(�6�|P0�hæ���� �ߡ�䖼oy��<��fq�h��/t^��0W�y��Nݿh`�&,Q4ԙ�����&�m������>�ȅ�-y��8�2 WC�R�t��L5_��Pã*�����Y'P�7f���@�3([w81W�������%�Ν,'#���
X1��7?��R��qN-�x�i��h��J65��sc����y�G�����U$,�<m����R��lC�{(.m���&���ԆA���Sb�����+�)��^�VT��ˀ�Q�n�>'	Ā;E�����8C���7��e�[V/����+L@�)���؆���W5�D;�ml�[1�v[Q�)�$�"���e��g�X�M��d�a����fwKQ�[�o��w�LBީ���
C�"��k�j8j��wi�ߧ�^G�pT�Z�O$���%e%�˖����
#6�7S+u�l?=U��z���!�Mj�8����v����35z�1Aީ��^�N��Mpq��1J�M�k�oܢ�SK�r���oS)k������J�y+t0��
X�(XDb��'T2��Ϫ��^�D���y̉���h��i92��4�����0��5hu�W\aMvk�~��V���ŧ᳒gF��]���!f��0�:���r�i}�l(z �Z���l9���u2[�ך�����m3��W�J#HU�5z�	��5Z�e��ш|k�v˂L�0�s���-�2��r����ZP5fe�3�)�ے,���� �7�>h�Xv\�>@[_�\@�5���خ�n��-A\:*�<a��|ʑi;2��1�CM�"���l�)�"�5�N�኏$1�jk'	{�Ü��O���$�[>�J�:��8Im7��	��� j��>�ۂmỉ��C�&y���,9�uIK.����dP�����%�ʜ@��r���fp���%��C4�.	b3au�,[^W�t5ȓ����2H�h����+��qͺ]�.�v�� �X
A��C��ZA��»���U�O7�b*Z|Zi'0n���g@~�4NeTW��*U��X�����X�1l�Ƹ���[9����۔h��iZ��Ŋ��#-��t�}Ln[`np���.��tʪ���@:�aѶ���A�ܠ�,"���p�v?K_]�h�?$̛��nyf��?;��XgL��)1������b��e8'�X�H�!k��/�e�b?���s�2S�戰�]8�U���۬�#�����m⮡PF'�6��qJ��)`_ٰ��̞/��1��VJ
b���ΠOM�iEo�xɅ����z;g��+ˏ>�u{�H�Z��}(_�;�`]͋X=����ߡ%6ss��01��o�ͯ5�4^��B����$*O�Ÿ��]e�zxi�!:��I����f��6�-Rʮ׿�Ulbo�$�+T�A��w��$�-���������ED~X0�n����q=e[�b@����(:t8� ��+g���5�͕s^^�c�^�C������_~�{k�]̡�(�I�F���>D-�K��H�[��lk� Ȅ�G�.�8�ڀT|,��A���m@�s��:��M��-0͟��g7�@�q�w��9"�"�$����~�~rm;��w%�3~��5��	�ȟEI���J@��;Du�{���-�)�ؐ/������?�ߴ,� ��[������P� �Cu�}h:ZJ�M'~CB5:�d���d
u�ӻ;�.�;�T��ŧj��&6;-�K�+p�0Vj��*��S<�����^�
�I+�!Tj5>Z��W澋O���^}�0���"t�j�>�)�O"?�zy nf/&X�[#5�����J���/�'i��Z��x�Efk��|@���U��v���P�l�":�Oa��|P�Nf��3��H�t3�Y���|ncS�"�2��	+��+���2e�EL�Xz ���9� "n�ځtl�����T�'Ǟ��P�x|"�J��w��s6/���w�Ϋ�+=q/����Z�u�g��\�>��fYlkOO9B/UHfo�y͜�8�Y����:��?sm0��ِj��޳=���%t�"��)	����$dӎ����Vȿ_>E�u��uN
�$K\�?!���쬓�s�ӡ@TC"&����CV�8�sy� ːpkdg��l���'�Ԩd��޹.�-!����@':�����wbA0꥟�o�d����_�
�	2Yl�_k�f�����������f�}��I���^�o��n�~�\+�5>d��$����"�|�j����ig�$�u]���?�Y@6r���Mf�t����O���{����!��<�IS�5p��K7G�4�ti��}M�|LL<$Sk�����	�R�X̝>�d�]����o�mP^3���q������� �����52�-�Om��Q�����[�5#�>(s���/	�
���hH�k�Y�2_�{A��RM6��5��w��ho]����D�C�P���MA����0j�}Ŧ�fB`����$82��Ř��[K�#� ��j�m�J�M8�7��D[���U��lP��7MV<C�.(a��`N��5��=do0�_yGS�:���]̩}�Ĩ��E�'�K��Ѽ���c,��B�
xS�~tzf��3�����!���f5�0�`B u��l�����_�JZy�}��!"�s��\�1n��Q����W.e�������%_}�v��8�3u������6��w��[P�7���z�s� R�o�o��U gא�{RӴ������e�Ww��#ĩ&��Q@?"kT������Z!��P�dl��r�y,�t��������*1����S�T��b�^Xb���D� ��[�p���y�'o�]����n�5�f�.�#y�a^5���;�s��a�����l�Xh���`I�g��q��1�T)���OZp�`�ia}֩���*��`Z��碶���-��I��gɥ�c1�]=)Pp+&tٚ�J	X������#�.9"�SW�
�1�f���sE��`WIrP<�/r�C�3D)Q��a�Ɠ�@��'�;��>n�\�z�2�m�SF|�$�v��s�TFL,k/8s��}yJӞ�e�Ut݇6rF�l���L8f�=��rR��T:�����/�$�E���!��/p�#Ŀ�gQ����b�'�s��,޴RmH�}�
��ێ;@�p}u���n8�`N�p#:W��6:�v�ɟ���]b���[��x�CjJ+?}�����a��5!	���X�v~>k��^�Y�76�Rۂ�={��/�yN�����*�Tۤ -� ������9~�8v�<������"!Y�H����%����YP�lߛ��L$��?�N�na�'+U��i�� ��w�ǐ-���R��}Ӌ�ߡ5�~O(~��y�Nk\�Q�,;�
>��% �YKy4F�N�5�%�H6l�d�B}�&��f�{���[#�7N��n}���#�h��r�;�mV~%;ѡ�jD��	<@e񙫾���\����Ҕ�����Q� �<ų:�����!2��Df�)�yE���Oק�sMY����8�:ó�Ş��}��sE*�������7� �vc"�Q�UO��$��Q�Z�r8��4��s��s�	0�#�M�̓e$\���P>�ӫ�;��i(>4DdӾ�����N�>��
o�0.�O��S�޽%��~6"~�q���1����� �ꙉM��M_t�H|8G�^!_Čs??`�������\n�2�m������ى�Y��c<��U��f����c֕V�<��i�Ph���v�)m�5ƫ��U��%���7*TA�Ea84��1��]oZ�s#�d��3{5��f�]��_��W�
��q�6�D]�ks_^��p"�ϩ�-Ӥ��	�.}K�ӴQ�:T����Z5o%��3&�AH�A=�<���r�5)�	�'Ɉ��zA�G^�J,~�J[��2ȳ�d 4`(^��*Q�h��jK�-�LO'�U�)���I6	A(�>�jG�1&��`OI-5=� ^te�����#�����y|D���~��{ʻ��M�l�4��x}���y���3 �D�8-|�WazWE)7@.�3����Ѩ{��ɋO�4��ʠK^�j�����>��C�@�f��`>�q�TK��|�:�̚�x��ω�����,�/�W&�i�f����al�f�3W���� ��f��f��H�S���t�V��Y��Z��%N�B�[g?�nA�P�^��������W�������U;kuɈ�Qޟ���_U��s�f�@��+~�\h��0 ���z�Y)J\!P��D�w������B��I�цZVpd_��e ���s]T3v�2���)FD L_�&�#�:���Ci��{J�ʣ���a�9G�E���D���5a���H�я#��1�F��G,j��,<7`���.�����PpE�Zb��Ѩ~K�:g.����Z^ 2�o�!-lBEsg� ��L��<%�-��ϑ�h�$Z��k�@$�V�K��`�N'�=2�R� ��_��S�*���CcO�q�U���LJ���A׆6���h����uu,r��(['_���i���y&�'Q[q6�(�Oy��Ɂk�-R# �ڤI���@�E㷆f�|��\G�B��>��LI�L:�؞t�u��=�}��P��K�N�8���Yf���$��<��/�V���gS��Q�h+:L�bi7�6S!#�"����m�
]SK�Q�����ʛB%h��m�ͺ����<JLg�f��dw֘S�0[$RY���t~���.1�=����1�x5Du嚔r-� ;���;��`��JIz�mؐ���n�[��[�0��R��"�V�-|c&�Q�$(ά�}�0\f�^��а:jY�T�z��>hhN42�Ǐ*�Ss��b��y��:��������b��R'�=�Oy�[���쩱 �oA4���:!1�l�����~GGPB�Џ�e�����F��� �]]�Է'{�v�*�Je��"4�o�9�~��$f�����=��:	j��nSAO6�j`����ڪ3�J�l/���D���1�"\{�5��-s�wXә�i���y��jl���rD�KS�TK��*����!�z��{���\�f2���p)2B.3�
�-��s�o�M�������������!2�;k��$\��{����B��]�k�P�%t|����B�=�Ƨh+���3�$(�,���������J��c��DDm�=(��(���E�"�����+��m*3�{Jr��"H��v�N拷p�o����H���L�����i�y�HZ��Z�U� �S��=f����s�3�Q.�z������&�Vz�������-:��-�V.)��Q��1��T�fgV쾺��Q��������N<����()z�ۜRc��	�O��09��;��'��,���T��y��T�r����"�ik���[���6z�U�oI�pMgl��xT'q�FP�+b0*�t�i�M��%)�2Ac\aD��`4W}լ��:>S�����h ��99�N�m�ꮫD4\�k�Ӑ�U�\�8d�4�?mi���)�`���5�9�����tJO�����a0!������T���h���SV�	�䝋�c~�S_�4�!ƨ����{��F �}��)7�c��9/ά�������>y~�
˄b��%; ui^�� �u0��G���E��؆�+ğ,m�� 3YZK�Wa�ܔ�gF�S!d7�RޠB��v�&xb�N�V~|����y8:����^�t.�/h`ڝf�P?��\d����S��;����>MU�R�����K~����jg�Q5�)X"��vq����e�;az��E�Ϩ�ΒNY��ި�.qz�-��ǌu���^5���e�_���ӯ:�ñ=*�q~Y�8�h,��wЋ�آ��v�Yb�,ܸ��~�"	��$����Rosj>�'�,)��"ͳP�Ok�ԓ��[}�T� _��i��wo���Ȓ�C)/�s��I���m�Xt#0��I�} �85�)�ĉ���'GD;:fo��ݘ�}�1�8��t/u��F�c��q:�.���Z��'H�XO�q*�$LaM*[w�;�,������"QH��Ј��J�/ʴ6�
^Z���cFS�Ǖ���%����d���8>t"ֆ>�6��Pw?[���&�tq��3��:����S���F���������+j� �=��(FR���%P�']Fq1��ٔ���|G%����x�UՀ5�M�a�3L�j�_p���s��_ٯ��I!S6��� IU\��.MuX�Z���އM�T(�eR�N�ٳa�<�3���`ܘ7Q'8;��Ch��$=~&�� {�`��瞒��YZK�Z��5��a��4<e������A��H�G�g���19���?��%��[��+�=g�� 1oLi��g�����vK�RG��W]_m���X�1���ʵ�đ�WN�������_;�贤�<'a����c�QQ�6nQ#����j���Q�-&���̚��1U9\�C���U�kU[V�ي�@����Bso�������H���A$/$��(���6P�]oi�}�Q���uU�^/�A�m��qΩo� �_#'/���n��E����]'L6�K������� (�9���Ƹ>{H.U���v���Pׂtó!�޲���Dsi:�RG��x�T�'��0
,7[z��ҽ��=f��Id4_gR�bB���U�K:�B�����g��?Kٕ�~Ά=�IS1�.�%<2=#Ǉ/�zVxu�H��Y�ZM[����_����������ղ��oim-����w��P�وP[��]�l�^K��D���Ri�Riے���)�#y���=&{�5��G��O�A�E��g	0��ްX
�K�ԑ�e�A�^��f��c�����q�`�1��H��^��&G��P �U�Ürz�(�˻�d/}bP*� .S���Z"O�M�ˠ�i�L�=�}UHO�ݴ"s�t���4C*��p ��<�G�G�� �.�t~��:h�L�D=.�k�_�i���������-��P��hjʃ�g��l�{�����47w�3O����K�������H́��?Ȉ��j$&
$aO���O�#Gա�s7ev�>\W�2k`(��J��Fy�c;�@ ԭ%��˃����qX���e/x����uk�=��n��{Rk��\Rsa���ēo@�	��h*s�=Y,���Ϧ�:h����Ij�����A�&�������'��XlxVHYEB    9620     d70k���>k��Θ!�:�H�0_��>��|^�w��2��j��%�{7&b�/���l�sH�0��ϚR���r��VN��w�h6J|�S����8����:W"��J�u������=� I��B����E�� �B����x�4���֚D�!b''�_���)G�2��e�A��͚(��^u�j�Hk���Nq3~��ό\�ƞ1+D�^���ޥc�+�15CL����߽a���IE�h�[K�Yk���<1�Cʪ�W�B�XK�Nxy��1v��5����������(,�����%]����A������{��Z+ZтMoQr�;�fZ�b�Q4%����C`7�Ca��?�5�
o_�Kz�TP���w�ɰ����x��)�� m���x(��ʨ��L���[��3	K=�V���^�l���X7�{��Zӧ�; �#�dĮn���%l�p�s�0i��^dk\�%�������`�|"��U���{v�X�O��hGL.�6@��B����F�@3��友��d<c\�3��r-�~����i�)���㐲��M���P�-�	�c�lG������#��������SU)kJ��YR�0Ϲ`W(;���{Bx&6�2��T�
G�bN&�4pY���Z%�Fd���|;�����UNv�z�v���p"K��VGg0=m~ʙ���~�Z.7� �/�J�ȗ���b[����T���>�FCs*#ޔ@��{��v��x�:���%qw��t]�q��q��;�����2�d�7>�޵�IvP^�1��\,�0A7n�w�!Xx��8�TP \t�oV��Y����)���w�r�)�9�'���Ȏ]�RV�pZ����[�]&-ؑ�U�����5��;I���G^�.�! MK��y\�~���y����fn﹙.��]^�i"���>^;�OG���(~LU/����]D���:�y�	�6ME�G g3�6b���9�z�٢Q�ƟC>�(+�ug�CU�4���*����o؝����+1��n��r��B��9�_^>���6>�Y�5G�y7�vk�M;m�q����}	ڴ*�e���b��_�i�!������B~���g�������@�ўP)�K48�'K�|X���oZ���>�ۙ��!t���9�B;f Bg��w:����|��']�с�/]7p�0  �dgt���+h|�] ���K����rVǾ�*��{��?�/�i��ʂ���n���P�.ڎmw����ܒ{��g�#Ĕ �:��ސ#x$�tVP�ÎO�}�my ��*���)VbvT����U�<;��.FU�a�P��t���P%lL��t`W��{=�����s���t��}����#���dz��>�.�o��7�(�~A���_�$�	#a�hN�Ҍ�^4y��-b�ܳ��҉m�7�Y�u Ɣ���L���܈��5�HiC�9�X��"7����ܲ:���TT�Y�Z�^�Ǌ�=2�qaΖe���0*M�f���.Z��A�H��e��駮߈ *�e��bH;~��<�s��}�a��dID�T�D~�����g,?�ͶnZ�������,��1d��]� M���O!I�}I�n0�"M��ײ��jg��B\�j�H�a�9��|_!��}
Jl�<`��T��ki�M�̸$�9ts�~�Ǻ�S�Y@٩�����	�=Qe�0lo����f��PՀ~�Qs{��'�� ���TuC��`���|�w{�ِJ��v�2���(Y4�N�aί��B�p_^�KUh����^&8
'4���5,�_�	@�vSA��.��F�(�ax������s����z7�Foݱ�#5�G	��7�I?|`��|��j_���&��ד=�u�>�,�j�
ϱlr�Y�6�b���g��7�01��>��ߨ�B��a�T��~Pc��/Z�w��`�-����MR�C�=_�|fnq��;�Q#ıN�f�f7V&ʩr]�F�j���~\��> IUYZ(bGy�ŭ<�b�����\������8���:(3���P�є��!�M�yj�bI�#�J�+%��5_R��
[�kl�RA�� �H���/������ʤ��N/�@V}�1k�ֈ�' �2��59�H�?퓷�Q3��U朴Ipc�K��O��|�[��\�h�M0�|l:�V��HS �xzl�U���&ǔpNT��O#�7 �Na��{�AmV��bE��Am�sg��3��9_�͟������c��m�f�����Gʫ�o�_q%�����K1I{b�L��0[���������Tn&��pc�gP-�qi7Έӟ�)�|��0U��ڜ!� ����-w���z�_D�_�,�ZGKMwp�1GU���:\J���"U��L�o�����d: )�*Z`�_�=<�1��Ǯ����
��nJ�/>�)6�����;pOLa32�<�)�:�Q���q{	O�mS�Lo	c*~LPr�g�ʾ	(]��œ�M���ͨ +�]�bц�e;��՝C�������ջ�ݔ$�ߴByN�6+����?��%�EL�F���{�v�s���l�����b�
�~Cg���:�g5#���8`	���|B��s���H�z�����Pd�d�q\PvDq�4=�����`RS�3O�Jvi��Z`ZS;O�k �K�¨�Xo�u�N��j��\�*v;(��4��O�=]���o�h%,5R�`<�bjX���*x�}����[T�4|''�%��
l��5:_Y`�B	�����@B�,�O�.s��~�'� `��"P�����y��s�	/*�=4���s �Q L8;ϯ�*�܌J�)���X|��/�qh�?ﯠ�_�w��X�FD���T��F���n���,.4�T2ڰ�.�� ǁ�GQ{&��LV�W�h�:����Dl��G���f��
��Jh\��eF�ɍ�ȫ#��?X/+����+2c��kA<���N���B-G�W�$�u���ph��;	�'���*,Y�������'��]��5�T���@�<��M
���r�bЁZ;����nUXw�l	�O�L>�SS Qf7��M�$�I�=��b�zM[����>�VVe�����U�v3I�)���&�����P��I��	Pԣ��.�׶����ˮVF~{�	���ڐQ�:?(H��j�
����1U9��5y�k��:$YN0���N�x�6���A��H|"�;�v��.Bf�'����_�.1���6��0����H�|M�v�a���t�3�����G��((m��H��z�����Gl���H�͟�0<�d%T-��q��q��fkl�?mPեj���s2ۅ���%��f