XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���\YmDze����Z�.��跅_k^8�����Ǭ�Z�Rv&v��*�M2~wyM_�X|�Z(FsuS�fI�8ZD�����璨:L�wu����pD~�Ƅ�Q�$�&>�/V,��A#�0'�@����㐶�z�gqĩ�:��$ W�1��pd�9"I�A%|���;֨A��$o0b�-�}��|�^�)q�7o�3:��?�3�}��h?�}m*��2��yF#��|�ڀ��[��i��J��P����K���������]xn3�����'�[����_b_'�T��!�)?��N�0�����a���P����h�a���?������Y+Y5SM��z�����2-��ϲT%��'a �LNi������x*�V��1L��XZ};�d�	�kT�uaKr�$���')����'k㤰�ձhOӳ,�G 2��ݍ�DWZ|�~�O*7��q��$��B�#a`��=X��Xq>����>K��g����x���dK�^ޅm㟸����k��y���hia- inF�; ��~�j;~&�9B���5L���-���R�#�,�]ճP&�����U`�t]�E�[��=`|�v�cT�V��Lbz $]�53�h�hi�3<D+G|Ϊ�vN=^��%j{8�_Q�cZ=��0?�SI�g�U�4K�Y�Yί�euϝ?�NI���iW�=�c�Qq.q>��g��U��.S�C�I�<
�qw�
�K2~H�:��g��N_6P�H1^l��K;}XlxVHYEB    6610    12d0��+�k�6�#' ��@��òx87��۝s�4���<�c�.U���i�[�*�D΃~���9�w&n��c�|?���8*S=�D)��kDQ��H��ܪ�c��
)���i�Hѷ�n�kB$����a�ԋd�%�f�h�Ab~f�u���cY���+w`����9& m������Gݶ�vDֲ�}Ju�^h�@5X�[ {���'�È�%�.檢$w��C���߰�w�X:�*��6���,�%3�ڟ6�%�[(��V��*sT���&�sIC�ۈ�/�v���\Lz���O�#e��Q�_��C%<kw���c��
��ֱB9�7���v96���tY-�#�-
�am���}�O�KJ�\c ���Yg���9{�u�+v��o��9�L�6��:�-y��C���R��Xc_�
=��Lӊ��_l�x�t�F�W�2�*9*b�O�7&�?�B�4�a�%��>M"k� ��lPɿ�f�h!���f�±�s�K�Fݱ��e)�([�t=+Ͳ����R��p�!0�p�5��n�E��lN����1D��@y�n��nǹ,��2`Dgrga��̸���=zoR�_�xzlDnL��U��U9�X@�R��+U���h�z��ȃ�~���O�P4�G��w�j/,��%6֚�g���p�E�<(\	}{�ɣ �C�n���U��$���s4��g�L���e�}o����D?�Z#ڊ���g�͇�$��Wr�kQ(����EX�0��9rz<��>���b%��敩sPZ�,���.M�Ь�~4�*�h�/#��z��=�����񿒫tg*C�Z��M�4F[����)�B�]�~��8��C���7�7��F6I�$��ނB&�{���I^��c?ۊ�I��d݌��!����f<�!^��u{T!�MߧW:*�Ve������ue�n�7U���۔*!6o��62�k��7�S����X�ks�)��6�]f���<��T;����y&]S��V@���%�%ߴڭ�;H>��E���t9jgh���V	O�̶U�*�@�����ٻ�\+�J��t�����\����3�ؔ�y=	�xb��L|��9(�y���ن��%>R���5w��~���su4>�9�����U���I�q	�p�5ew�<	�o� %�*��~`�a(�z9�,ڊ/Ӡc*�+��o�5���κУ���[�]pY�X^VP<Oق�d~a�v�i%p�g� 8��@m��al�>�ڠG.�F��ۂ��\�o�ގjP'�=���\�#7>K��g���w��qZ`N��)>�����ۭe�;�����<%��1>��e�׷|}Ѣ}��?�&��O�n=s׫yq2¼"��L�VÀX�gU:MB ~l���/����ҳ���0&�{�.$o��Ǹ�^���:����O"���'��n��"�E�V�{M�)�f��؞���lӇ2����!��T�&��YgP�^J$L����P�}��[�y"�]_�#T9aY���B>v�Ψ@.�4��[e*7
P�K�������<7ja��s�Z�!����+�;E�~_J�P1��|f|��]x� �Xx~a���� ����>�`!�t7X"�ΫN=����M��֧7���G��C�&���u����Pi�l�	�F�I��O�*M�����E��������R&T�i�_rhwڣb��&�Ac�J�lZ���	i�Z�}�����ū�m:K�I냢���s||�?�u$ ��P���	���Xf�<h�7-�M���+\(�[�$�Z��I��To� D"���%S)�7��:��c�Ty3w ؃�g���ϩ�5����.#�@$Fě�í��'T���-�H8�ѫ�>��~4�[���je�Ut}e�.˄�//i�e�8���5�]�QWb�]
��r尌>�Mx�����/���W����~�]բ�hFQE���	#3]�NX���V��W�I��JզXj��BC|Ƅ"�� ~<��&Y��l�2��H�Ul���Y��a�p�ɳgy!k|�;��^6|�<>�']�l�\��归ܰ>k�����v^�|�	# J1G_�����DC�^Rjn��ބ�*\���Mp8�Nx�Mʨ$����O���$������ _Ol's#Hl�-�
;�0�ۨ�]-�g������Q��|� ���Ip`��*�Z�_���x�WU��R �O���62}�ˋ�4�I=�za�CX�?�`V%��bn�{6�`f+�v�W>�fw��6#��`������Ů����%�ִ$"cz�rPd���T�z�����=#�.�^=c�'�H%���1.`^�� .�(�m����~����=���uIX
�/b��\��(��Ѿ�>������r	0N���A2� ��kJ �����{���i��@×h���Ǯ]��9��H{�(o�*/������9���P�0�2��1��\P#�U�9�'������@7����r�к6�b"�?�1��lh�P��{3�Қ���A@��$�\�/��F�s��b�o�Ƙ|[���BY��*je�jZK�����;�WD�۵Ju{ i��"%΅Q�'����V,��a�T~"QA��48W���j�-^k���>���Uϕ��=1I�*�S 6�m+�6�P<���4����V���k�� V���,Թ3�~J�ʟ[`��7 T���D*���xN�˾a��;�N^љ�09f<0&,�_�����Q�E$:@������s����>z?4��
�H\4�=�z�P�$�y����ъz�w��Y����t��|���
:�����h�@���x�#�ߚEc�
�9���焻0ɾ@�q7e���\oSC�<X�F�?W��Kl�R%X�ᐴbW?L`B/�s�|~�w���Z����3VoN\P�@y ���a��sd���O���/��#�Yذ��8��k�>1]/Z�9U�d�h�ƌ5���e�R��?�I8R�gn=��`��O��9� �����]?u��~��(S'k�� N�.�r{u^�х�;�Aaк�5-�5�����ƣ���P�,$��r�*�������	��7��m
~���+Up�>�]���]c0���]V�u	�i�Ӭ�g��9&I��e�^���K�R(���O_p@~�=�����K�B��L�p�d�*Wh�od���v6��X%���R9��n{�k�U�?��Dmf��y2�ER��S���Z���ȭ~�V�ƙ\6��> ��Ð��L�d���0�ݛ;
}�>l���\���jڃl�D�|�K�#@Ͳ�Bt���{������>�dl4����]��aJ�͋�ܫ?K+���k�]��e�k�ɓ���S��l�XX��c`>���ړ���-����p�H�S�.����.�p8(l��Z��-D�D֨�#��DP��L��i-s�B��R�3���:k��0�B7.%I2��-
�6��mM��-��7DLXE0��h�@��Db;Q�]�N�hrj����`F*�����/Y��'��R3XXsR�YK��a�����m4��3z<\w��cbl����5��8����F[V\�=CiK��g��^i��S�9����hT��v��6 �����(���w�}l��5Kd���4�O��}�Kt
�}��0�V�B����"Btce�U�)�O��%�����I�*��~1qQs�%�� 0fL�b<���V�y�OEs2%c���O�
b�N~�AG,ǫ�e<	PM�,x��-��?�)��\=\-ޚ+��!��P"]�2��q��#��(� �������8��>�|���J�:�	˓fO�2%0������#J��D{G2���wܺc� �jy�@�� 9:�cvɗ��2�m<Q����*��#o��R�����&#�0���ߗ�~V����Bb�E7�'�M���Q�9&������7����������@Tf���pbH���;�Յ��D����ιw�jOa��� $L=��L�p���z��6 /.sx���5�Lktu�|��2��y�'\�w	O��=	_�A�Y�^�:1�؟�@,�7�$�N��[O��AG��"��*�0��_	����2����q�!����a	�b���w�->s|�����&�����/b��J�dՁ����d@�^Tx�9к��e����:�U�-�ȇ�.eg%��v��|�&���7�=����P6��hH]�at�\ z�"�-X,#��OO�R��1���� ��)�����3��ՙW=#7��1k�PlZW�ri-@��5��I�FЌB�߅T@AR�{7݂4���ّ�H������M#�)q��bW�^٬W���H�c�>���~��=�������ã4���#��XF��M�����x%H���!���v��nRb��i����I�@�쿴\a���2i�7���=�<ǔ��$ud�%�V��<g��0���#�Pz�:�"�|�7�2DaA&w�<	���%%��Z��MAJ�|G�>��o���$]կϟ������t���*�򲩢U�Qj�e�ER���T�Z�!I�Y�K��(}ow��W�~�Ġo��]��7���H9>�t;X���6��W�Sͭ����]�!�J�X)Mָ���T���3�����{�e���e�~���k�������9���?sdU���3����Ew:g���4�8	ɠ����ˁJn9�1 ����Q�<	���71g�ɪܣ�F��Ri�J�Y.��Q��`