XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���0Ҏ�W&=�p�(��k$�c`àXq,�1
kN�n-&�����R8ǰ��8Fm,]��-TH�X����X"�t�x7ߩF�D�|��W͐wa��rC��˱e�7\dC�]�L��Joq��!�� �r�A ��J�vjQ���Mez��Y��(o8bԥ�LI� L�>��nO��b�s���� ����;o��B���"����T�6£#�����"��%��ݾ��z!:�c��.^�@AOE8�Y�Ni�߽�'0�N�WS���Ll�*��+M�Ъ�j�-��V��W�/�SQ<m��㙂�kE�O:5�;ܑa�� ���`�dT_���y����c&hLF(L��;!�3,{驝c��bϻB_��I~w�'Z��ף�l"���
ދ�	���%�{s�z�ɩ@�j��gSy���b�$]��bJۂ��6��!��ߐu#�fl��4x�b�Coh��G��`�4>�a?�O���
��M.�n��G �:���cε�,�'�2#p���FpQ��W ��R.� z��3�\��5�t��!�"�Iٰi��K��m�7�+�>���e���i�s@�~7�����}9��J�4�����7ƛ��GB��c=?�R~o��le����M�SᩕL_r1y���tI��2�Ҫ�g��!�d���;ŊD��T2~��Z\�k�(ɡ�O�1?Ƿې"��d3���m�U�_�<C�j[��ۣ���w�bH�`G.�Jl1��m\�kbu���\��Z���W�>r��XlxVHYEB    aa52    13d0�U�E�꧛���Ƈ�T�٘9[E�6@~�Ţ000����X���C�Y�^P#��rd���U��5���PV1���V�b&��,�K�@	�2��a�|fP���6,���� V)@��3Z> �z�+��ϯ��Ҡ/r�܄�2�wGOaf?(=8��c�s��w�`%7���5R�F�a�Bg�^�Cw=����U�#]K���(�`���n�oe�>.��s����d�ī~D�- ���!3T	T��0põa�M1	�����5R���L|z�ňգ���n�O7#|���l)�HS�\O��/ea" �ý�5�4ė����Ǩ�/������Q�HovM?�bA���@8�T��r#���މ�.�H���M�Km`XDE��7� oU����6���Ց��%L#�d��U!�X�k6��Rޡ9����H�A��T��?��US�Y[s#7��"��ӕ�.Z�_fo���z�i�9o/v��tn�8�KݗW��K���ֹ{�s��%n���=yYz$��wz��8d���kj6`�M洫�OK��)��Irm����d�w�+[p{��֩�!�[��|���B�(̪�>�� �W�4���9`.�8z����&!�~!����{�ovk�7 	�^�!<��I��k}D�'��)f��p�X��Fj(�h�	1�����%7�bQ,�s`,pQ��Ba��S4����;��8�j1�`�嘡B-�S��J����%U�@�"V.�Qc���tr��zme���E��8M%��a�6]�Rc�2m�%K�L\\��Q�2��a��}�II^k���55��3�9~]t��l�;Y�:3���,���"��t�j���o�ǯ�jؔw�:��C��&8�{���O�ail�s�`�a���Ev��v-ve�%�����i[�C.`�mY!�'8�b��}张�|�S�3p��(�d>&��rT�y���wb:�R�Rw&������i�V���)S̗?���]4�2E�b���������S/�vɱ��9�z��~�!�cz� � �J������|΄*�ۼ��1��2�~[��pt�[Y���S�h�)^��9X��A�N�똑���ZH-e��<<�C�c1��i�e������\ �c�6�J�/B8�z��0���]=T����^�C���ŝf�h��[��j�T\+�7����2�O�?�c}���*��R��T+$�n�G�RG\���8�\�
 n|aژ��=,*Ψ�/H���y��' ���L���w�@�Xu�t�}�
�/�&��
?%
媎��J6�{ga�`#����2��+�Ea飚(º ���d����C���4SԚ=�vv]�c��ύ�aO��p48C�7����5��Z&|���������3yd�1�{&���h�dl�ADK�:�r�G�������'zqL� 5��9��Z��������6�@]u�SAopr��lE2����\���a�Q�>\}�^>�F��qB������~N�� �#~����צ�k��U�e>�e%La��;����;L�1�W���lZr�D�p�0}�e�
;�����C���뒲.$�:`�Gt����m��:�GJ�6,
�|����֠�Nu�"��p}�/��h-��Im��֓1�pV%V���-��sO:.��+]'~a��~�DT�������/=��.׮����L컫���}j�o=��h��߁��x'��dq���$lkԏ�-�����ƞ����7Ș����$�cͶ��)>K[3��#�IEI���q[5N���*s�q�4�6!���:
�vQ�W�]��ۓ��8�
�5	H"��[�n�pW��`y�S}ޜ�����YJ�ḱ�u��,LW��
�J���ѱU�Dn�bX����=.�z0�i��Vӝ��j�j�Y��oմ۷Mx��ߒ��o�cO^�ݔ�fM��3��r�i-�ech>�`L\0JhsI�`�WM�&���S!�\�33���r'��㳻�[g�ǹ��L.8Ua:K|�y����4����O� ��6��;5�u'�ːDBYC���h�`0m�~�/�t"��{�8�az6��NV��<��qݿ�+ٷ_'|�7rO�AH���0�p���F�4Dפ�D t�ym�R�W�W�l��l�8s4�[pW�{�`/r�r�����슴^�W�Z-V#��۝���ϳ��=�������f%�95p >�ŉ%%;�4O�Z�����A���3!99ɴ.�P�Ef��-1߭U��!�ؐq'�}��U�ʚ_����E���՗ƦZ�����w4�c:��~��VC�͛ݻ�?.cd*�}�����?E�ז&G�H���\�E�wO�Z��+�#�H��
�UtJk�������;�4�������[�ϐu"N��QF:T�5طj'�Ƕ�_0�������U��$��6�m�ٌC.El3��3^��(v[i/���z���G��G��|"eU��_�,���8�(�W0+�2�a�����r]=�_��*�s���4��*Ҥb�t��T���^��p �!^�����y.&���e��W˪�и0JNU!�CDm��E�;+�m����#�D��J�ÁHϠ0���՟�N���X+Р&��5f-��2��;Qi�xr�tX�]j�p�	2�N�[����٥�a�yƂ��� �?�?\�Ry=�@��m��Ҳ)�at�!qKu��\����v��0���M��r�k/��bO�Ct�dh.nC�j�U�)Oe�>	�pF��t4ɞ�½U5��>��_
�X���}R�����]������=#��v`�]��-n�i�z)'�֯��4P_�@�~�/u$�Boz#����l���&�8��Ԛt��xLr}�41��e���v�G��)��v�u: l�c/�*]KO�r��ŭo��șHv=z����Mn�}���78�o�qZ�m���^��>������;f��݇d�6a��H��`��yd�%VAɔ��8�|t���jw\�݌?��?��������/�@��~�9󦻈;�t�D�|�ǮY/6��b�5M�Jh+%����s�p�+r�G��<��i�1����ZD��R��������X=O��Vg�.�i�T�y�0�U�G.�zӜ�}�ՙ��儧v�|r��vA����/�X��c֎�i��~���������\��#~/��b�j�}	tǦ���r��Ќ��8��R	��w���,�ImT ��C1�����@�!��.�%�")�m��q�{�
��Rb���I���Z�h�gY�ܖ\O!8u([��a]�-�����Q���g��6�o�շx�Ӧ�q��U?�s=�E=�F^y��å��=�)�N��ş	p6j=�ZM�{���,�s�WGy��f�H��rB�N
,Q��E��|'��.h,�iR���	>�mb�B�AD-�?5#/SV�޾���a�NCMG&�{�eUΚ`�l��`�G�h�N����t�U!��� ����
ݷ������� �k�T���7�7����Tx�O��_�i.�o�9�i��ϱ��i2D��W���ݠ-䟳�K	Z��7�e_i���Qd�6pkJH�~uu�eGN�G�]v���$��ݾt*�L�� 0�r���>|]��0��)��%�Xoumv�����Լ���u�4�����vX���:��/X
��~׃�X�Xx�m7��!����<(�S�"���H�WDq�w�|���T�a2�����d���r"؟ȏ�A��@d �������9���E޴�"�������4��Y�'u���� b��R�d����DE����/�͌Qy�2À����_#���qZX�R���>����T�R�� &h�C(,Kz=P�� 9^S���2���x �na���)P�rʸ>�3�3$�9��<x��^)E��m��JŦ$Li8�����W`mE|(�c[�\�2�ut�6s)Ʉ�����;�ND,�n�#i��rQv����Z����i����y)lLR���~�0n����O~��߂H��u~r^��^�s^���"�Rͤ+�=*�V�8ϯ��Z�UbTL7��.��D������ޘ�k��cL�aܘ�ॆgU��Tפ]��c7���MH��׮�X�^�FI4r�����qu�xq��P	�k~�$���F�>��������r֍ ��K2v�V3x�!�4��V��p�4�����y቏�0�"$R/��H�g�(r�����6Ch�&��0r��6*�S�x�~t���w��g5�e)D�fEL3�,�qqAp�%�5H �<S*�'gL֭���x�r�5�M}D�uF�>�v�z3��#�Xdc�Mk���������X�m`JWsw3j\0 �'��FMr�BG����eG.�n�<]!׳?��4rO�kJ�����b#]�֪�G�(d��k=��s���|�0U�Ӡ͠7?�u�wLʯ'0B�-k͹{8��_�n'��U&�zז�LM^i�zQ��@qek��X�v
���b�_�Fw	@��L�ѱw�T����h�0��Cճ֟V��sK:-Y�"�?�Zbҩ:�@��$����*6��9��a>�M�y,��/'�FBz��ĭh�%��(��E[_as�9���S�M%���8���n�Ӯ�E	���j�]�� �,צwfӣ�F���wC8���L��t�'LP���<hs�hE#�V!f&�����M�"�x��N5�Ҽ�J-�&���ɱ�D�~�=µD��JeM���ص�0�Ҙ&Ї #]�P�kT2o�yܺ�\d�g����Ve�s��-*�'�,��$b �B�����������&oi�p&��KJ��;d!���������=��V&R`ʟY��1�-���Q�ǽ|pǏ�r�k��A��ɱkI�\�nBr�:Q
���Ʉ{��,e���2t�[N��!h�{|BB鞟0*T\<|L��(w