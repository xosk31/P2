XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���"��=��Ù�ޢ��l�X@,���N*�u|B��1i� �F���J,����0��Fu �}��U����TK���_���`�e�)G��[�?=+j�6&^� p����ݠ������z�6�w�t�j���t����(� �u?͓�<��S�7��ee�ɿ���:��2�͒��2�8J�He��awyT6��yjW��t��������P���KϘN9Y�N1�,	Z���q3�� ��81"���^p������٬���P�	5[�f 	Hy�r� 9�d|����&'wj�]i!�2�K>^��#��u�ɹa���9�<{Dh��2䂟,��'�-�Ё�Z��_p7�*3䉒F�$��mm]�J'��q��Z��r��`BC��O^�k�~U
ต��mO�����^2���,,�Ȟ��}�����Cw�(��&P�@Wˈ&2�O[*[�8��78Cg��A�;�^q3�}!,������_YD�~9�^�m�B��i�d�H)��_�W.�:5�� �u�ո��Bɼ�t��­��6"��"T�%���[i;�^1��ޡE0�9�ho�rs4�=�KR�M��wv�@����-�ͽiC�5�"(�(�.R2D�e����DAe[�B�0�����S"�1��H��_�;��3���0=��_y=���/s֡7P��M<�4��Ǵ�n��6���P(��c&w�����4�Y%E$�H��w���N~���r��jXlxVHYEB    3b6c     e50���{Cm������n!§�iw�<꼉&J������޽�&�'�%	x�^��%��=F���ך���f=('6U ԏMI~�**�	x��\@o�����e�x�Y��ҥ"�O��P��V3,ѩ&
���ҎT�8�����<�v-�����7'�TYlE�JTР��<�u}rz�_������E�p�uِ� |��U�jF?��,#J�5*�
�U*if�0�LlC�D1�7����A(��| ������\�3����UY�5�	g���ٴW�@e�Z-!�{{�(+z����,Eׅ�苃Y�]���B��[��h�9����-HilEsDN���C`=R#I��$Ei��n�31�*w�G�d��3�3z��P7�HM)���.}�4
��Nro�7eŋ��.đ�E��&��0h���ڽȣ�\�p�^�Iע^"���{������{��ɽr�(Ç����4OM��ѐ�n�3��#Ȕ0�~��5f��w���I��Y�GC-���uE�n�\���S����J���[XK���/챷#V��G�0�w.�a3�Xc��Q8f���a�<,*!U���c�e�J-_~�;���	�y��U@���<����C��ҙ�y2І���'���Y���C�?���H
~�3Έ)�����n��Yx�'��&�HF9�i����M�{�k��,�l�<�<.����:+Ѵ�F�y;@ ��8˳�{(Zu�k�P	��W�GMs�U*���h�`�8Fހr�m]|��9�+����7���V1xD-���p��cw�ёe*3��8z�0w�F�N������7M����`)"���^�e�����*ˣ;Ȣ�q5D_�#�g���7[�&�������y��kz���4}�1��3�Vu�w)�D�����⽆Ga��	��s�����˺e�[53})�����J��B�
;�p��{$VeG�񲺭�~��tq�X-PJ�A	J5Jܧ:��6�EȄ�j��fJ�-�0��(�#��PWU�T"��e'��OC6��}��}l;5OR\%���e
[�w7_��@XŰ�-7T�_��a�ýI7���r�;n�1� t[c�e�g�z��w�#�{�pq��Ͳ�/�ĝ&��O1Ub�>��S=� n�m�9�-Ŵ�-[�dqi�C���U�Hߴ�m�`b���#���&O���j�O�0y#�`[�k�����t"ڀ}6�m���a��'�2�>��xP���s%˽]$Z�>۶�r*�H=�T�r�o;��[*�yWm�V�8��j�g<�lJ�(�yq��K�k�{(��q׍B���\C�1:F9o�D/���bU���e~���U���wj��k�\����NT�:_cǍe��T�$�_�������Ľ:͊�9}Y��k$�'��VIiˡ�|l-��C�����,�

������4���%�;Kz���ިA��^���T�y6��h������g�2�_�q��(��Ŏ�U��:1V��+W�~��bo��z<PF�(9e�bL��e�/��`i]���?�`����?^�x��]�/"�8�,`�x�� ƃ��Da���mO�T�¡�\�-
�j���fnf�R7���Җ\��@
��+9�<����Q�>�!�b��r���%9Ep�_�U4�_�� i�%5��a��N
�CC��(���r� ���L����e6H�=���Z{i\�֞�o������0]G ����ߙV�"�Z�ȗ)�'@_����
��ݾ�l�{%�j�E�.��9��t�93�~L�����v4.<v��lc�#�Β� ��zo������K,��.�)X�ld��~u��8yK��3� �玁�2r̳�:�|��������6ʠ
��$L�H�gR���������d�-w$�����:٦5���N��D�]��l���Z�߼h�_�)99@��c���q��a0���Z���%�)���sh�4�� ��B��I�]���AQ�HԎPL�3�\�d�V��4��2_15��s�To���$�n��9���U�\~:��j��z��-���4bɖH�C���h��vt��q)��%m���Ћ�y��༃��˭�}��t�N�kR�G�@嵟Y+zdFԙx�Ъpc�n`��D�aG�҆e��n@.Geψ�J�r<ݿ�����]&z��L˾"N �.��ι��Q���C�I��2l9���!�����<�.���< 
h���90=��ռ�����+�j�	V�w#��|���D�e�������H���\������?�����n0-H��X����ֶ��:`�T�v��bh'A��k��?��贐d�t���4n��~4�����3|6$��hL�F�`ΰ�y��膵0��}Q^x���U����`S�Ƭ ��V&�s�+����E0pDӨ�k:,��UU?7.�����ҵ^�g��,Pzxb�eÚ?�֊�(�S�eL�l��v�xI�����.t+�C����v=
�� �$�rM��\5~\_ D�������"��m$��	��CE� >	�P�K��W�5F�л��r�<�ϼ�ݏ��,����\+���Z磔���G��+��y%܎��!��ʌ3��S�]�Qݺ&�>�X(�i4�4J8�WBpo�:��<����w`��V�J~�� X�rM���1H��P�U���,�p~�{<������61��|"aD'��	�o��THЕD=�p�����6T���� �?T^�ex��L(�$������l��zD��cyOh�a��m#Lj��7�j�}��dW�YӰ�f� �X+��Gb=��oBb_"�ꂦ�z�rD!u^���OU)���ҹ if����{�ۍ �ʍ��#�*�@@(��a̗��ȑf�+ZJm![�g8M.�z��=��[�=F�o'�����߮O �4��nD��<��H��*�~�:!�s����Yt��#:C���Z���o&�lU_�6����������4����Ai/܌��ykM���\�H��m���~u$l'g�PK�>�;m�w��y��H�N�cy?��!�N�>�DJٗ������M���<�����ڽ��J8x�s������х�`��pa���A�GB���o_��1K��$i��[I����vN��o}�'KCV,3�T��}�|�~�B�	)� �H.�d2�	����}`.�P���c?	%	Hs ��t� ��#��'-E��WȗC� wE�v3�a�6pL�6	�o�p���V
ɭs�6�}<E�����-�Q�I��ˀ*$��/�p�j>����I1�f�(Fh�̘H*��O8N�?24$�w�2F���<���:~:K��獻�6]�DA�-��Y����^,���ւ�k�=|����Y� Ǳ��U]�#/�5{����uVg�A3/�~����9�W�Vu��M�1������~lv̭6����P�8�11�!F����ٯhpF�hԎQ���@�5F�8����JF&�yߌZ�� �>�usL��?��a�ꪳl��j��K�0�D*,��T�WE��j��A��ʠl�j��!���9BYp��AM�l�����Ģ�}@��