XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���c�����|��w r�PQz���+����H�� ����!�E��2�3���H��3�:�$݉*��1	YOVFD3��12�Hf��Ļ] <J�S5�+񛞡]x �xv�ĉn����jv:�n4 �sd%{P��r�+��Y͏˘r�E؞���'Z!/�Xx�wD�r��,���B_���vWU��{W�|���b��٫c�k+ϧ5~�-:[_B�d���yӂ��H������6��̲v��0�_�z��lkn��qZ�P�_����m�%�*(����u��5��?S+�@*Vg�ﻮL�VՏ�����^Zё����0Oݦ����0ӳy�<����2(��v|Y��`A�Dӑ��f��#R�����`�@s��>�c��MN�e���#���Ҥ����{l� ���.��Y몰�=C4�:���`�c��j�:z=q�s庂!�ڨ@������y���o��u,�/��IM�2Fq7��l��P�nͦ$���q����?���>/?�]����X���'���E<�Ӧ<Na�H��\c���k�h�Δi&l��К�9k�}8�h���Gp�w�C�ل����e�"@o�\}�ޫ=I�Rd`>�E/uQ@��Zmyod�����d�E�(�/9��9Yj���w��:�F�?2ql���/xm�Ă�R�>���r�O��jQ$q�yPޏ����cK�6��+>�>|�R&/��WQ�:��'��#�Al�I88����%�$|>��,g�;��8pXlxVHYEB    2533     b00�'Ât��E�c��P�l�ɩ_�`��?�to;�Q��a*<ܡ�uǞ�j�:2(���dW�P��',>@w�o�ϧ���4w�H����4���~���$%i�S�D�ev/u�'���p�\��} �1��S�W:������w���O=C��E�������CSll�jB���]<&�i���>L�<�����M�g��Y��<D��ύ$���U���dS�:T���X��So<����}�HL�D\@c2�wu)���EME"e3��c�8�F��ɑ�:۴��M�����~������{p�+I3H��:
�6���)Af��������j��^Č!������(��d��kuzS`��	 �o�{���qo�����ϙ��$'�����i�����/�Z*u���b����u�� ���[��F!J}�P'"6�v1���1�ua�� �,C��1T�����˯�B�����R�4.�d�AjL[�o��q8�w��s���G�K e��J�����MR$3��XG�k?Ե4
V����ҿ�}
�>�B�Oo�}9�[��t��^x�r$�
z�m�p��:CR9��Q���쫝mMT5�{|К3����p6��R�ꢧ�\�cqd���G�묏��ua�5��/�/q&�Ԓ�]*�_2�Zg��u� YLP���c�'�n�����h�������e�_�����,�����b��dl�{��)9BAzkY'�;ȯ�:ES��Œ����Q%v�-�b�|�5�C{7:6A:i��)��������\� ���z �|n����$�;�7��ca+?*���z�jӦ�0��>���B�c�R���u��&��]C�������O�aD�7`��"��P=H�g#��YDO����C]Ah�^P.j�=�w���0r�ў,�g��Ҝ.:��o�B�RS�ve�U�2[��ԣ�-�5Y���c� ���J����/��u�����y�&$x�.��?�����Ӿ���݃1L;z�k!�[��������r�)רr� &�oGC��Y��9uRB9������XJ쯃EC�w��	����E� [b��i����ZMmrϏy�� �M�� ��߻Dq?�L�F���m��ePCb��d	�y��E՜�"�Қ�����Iz��?g��]5F����$DOy���R�Qm��9!�ϛNc�G�����F3��/��A%�F�,_,\��w���㎰$8q31d^}�c0*]��?�c/�=�(�����^���2�r��W�W�z$�����$�-��+����c���f����+M������1Z	ٟ��Y���|�6W����U#��i>o��j�~$�b������_D��ۭ��>�:�k\����7�;Z��N�:�`�����pMQ��a�`N�׏W&ji�I����mzN��:%o�+�m#ʵo�t�d󆟷�����=� �d'v�&�HC2!Hop�CPm�	��1�tl>�2����+��DF�ڙ'�f�HA�]]�\�����Ԏ��N���݇L�9M�;N�hk���ȼ���������7��l���g�i���k���]^�����C3L����7����9�UC�s��'��p�K=׺�a�U:������y��^��0+�����#H�V��~J��Х�^�~�₢�L��������
����ʅK� ������%�� ���uӻ� ����� @ىt�/���@�WQ�ջ���"ۡ_r�b>��e�g��( ��˹`:˫h^��p%|.����t%�R�l��Jڢ�pp�m�H���_g�E/���Q;(�]iư��~F���2>нZ�f�肿��9�;��0�1�j��_�>�hP�⇄=c�Y�H,u������i<��T�LW�Q�C񯎏��	ɫ:s��qf�t1�n"sM��о�8�'�>�B8i@}=3H?�ndE���������Z�K�V�@���A�P�����4�>����l]��MQi�F����2��
��w�a��g���M)��5�1�U��c�\#�.Lލ�W��kH/�j��?�r, +�Y.�)B��o����L��x\����C&O��5���>�4"��;���e�km7k�]����G�q�ՙ����~�y\��%����_��|oMGH-Z�9x�F T����u{f gv��C��5{��j���C�����V;E�|'���b�>���ՠu,�Ka��q��#�w}J��l�_�T;��&ߑ�<y��<�.X�g	�3W����8t��G���	Ԭ�C�`�ȯX�F�F͠���c|�%�R� ���������+�]|{g�|�`$:�P�ނ8��ҙ&$���6�;}�a��Z<R�����"��M�yL�r�~e�w2qg~�`7SK�&1�djJQ �uc~�6�n�b�C��3��V�mi"�VR��gZ��"(Y�)7ڣ������h+����H:�̱>��C&�w{�<���ŏ�(]��O)�]���b�v+#h�9��R�˴VV��ݧ#tAJ�����������3����'�`�ԧS����{�^���Uҩ{ܕI��[mv8�p�T
�#*��\3�<.��7��)~}���!�6,�W��+�1�����n�Lۍ���ty�@��i��*�7��I�蒅!/�b6%���Ʌޓm.���z�zO6�y����z����6P�"ڂr�+�u�
V�A�dh{i��"Fn��<$s�8i��*��5�p"S�=t��