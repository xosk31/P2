XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���4�o�8�,{04}U���5��
veUg��-���c�Y���.��]�����P;0V�`@i����~�D�H��+ȅ)h��W����%ܩ��E�0�wt��5A�}�!�![���	���6o��-��dd�n�pǡ��R�̙��]����C���f��_�m�;��A\!y2�v
ǣ���ͥ�����ú���Fv����y���^�%i�jy����Ma�f��1 3*n��[�
4������W")'+i
����z���m�3[6�;�x�Ā#��a����\A����-E��צ�b��z	O�|8�2koAN�=eS����,� ��[Z,����]F�� P=���}���3�(��y��P�	B�,@�PK/G��<�6o��J8�����fM1%�� k	���p�Y��(*n!�-I�Ó�+�l���R<�o2���Y5#���@�\ZH?�"M՗�y���T��O��_#>CX��,ٛ'MK��a\�iA���[�[�eY|���A<b	��j��l!S�σ��#b��S��nkؘ|_-����/��z 7�1A�NC���+bH͍��̍��I$;>eT�[<�ۚ�y�ν�KG5��5)<.=����9P��]6�NO���&vՅ�1RL���}�6\�e���d3��x.��1��/Ju��: �����bT9[��PgP7R��3o��q�J�=�6��;v"��;H��� ��e1v��k3���qs�q2�" s�>c�,�NfbM9x�WXlxVHYEB    15c9     850F0'�-�ZM����Ƣ�g+M��6b[C��ؕ�p�fֿ[�
A1�L33p�M�.�{��
��� @b9�	B|�?q���|�dj� � ��PZ$f}`�^W����v	�7������z��.�.�c&��4��aH�ţ���
���4	H�G<���uRD���� ���!}j��5���_��s�n��BP���_ɚ�{�T�\���{M�V�Ã&�,�c9쬼rg���G�m�#ii����.�d��R�w�ٰ�\�_#UN�0R4�b��c;ԇ���߽�#��`��T7�?]�K}a�̎�H���*��]�C岞�~�f8^�}.�m 2�+�� �0�)�(#D��1Ӡ�1LohxI�/S�C�Z�K(6*߬��	8��V�:��b$���?K�&��G>;��Ú���'���\A�M��[�Ծ�b%��Ʃ���ޣM�BC)&�G�Jրv9y�)�qc�G�<�ϊ�?8�Mt��5娒�t��w$�����Mo�?mf}���ror�q֐��׃�@\'��B�[�Ȱ7�'�z8�#˱ƨ�b�[�6=k����V�R\���:��KO��e�h���R`�F}�P�&0���r�����c��3z	m���@�nFW#��\�F�1%4��/�d�h��=*D����
��m�$L�}%e�)��]��}8R���E�����h`��(�7`����2�V�����i��.�r$fd�B�u�p��}���b~ϝ�{��W x4�н޿?I��6��I��(b�w��H~�g��_�X�q�I�����Pd+Q[��Guչ�l`��ٹ��{_�m�����)��q$��p�g�p!�n%�C C�0�E!Ͼ�e�Dl�D�~ :hRlR��x�\TwTDL�50}O�'>P�C���&�RG���0�/!�$V�ҝLv��N����uL]�b:�mHH+��{׻'8��*�����V\�h��0���;- O�-C�{:c;�A�s�����?F�s��t�c�NJ�uX��Ǽv}I%��q�Ň}J}����g�8��-�~�ˎ3d$M�eŝ���|�-;M���4���������JG7�M���X]^�TӊK�.G|�Oh��Hb9��z�Y�x�>�C;	6F|K�h�.gX��R�i��b،�'B�0�/Aˬ~tF�����L�$�z���y�f�DP�҅Z����{�5n�^Q$KO�k�c��+-����/�(��B����d8p���9�Jb��H��=a�3�J���q�@��anh�e��cl?����ߧl���T�y�Ɔ�^��L^��=@��o�w���yU��ə�I�O$}�Bw�.;|>ѠR������A�j�<�Ve⎹i��Ã��W�H�'�Γߞ|�ʿ�@}_�+�_qZ�>% ��ߑ�o�5�a%nw+�zׂ\�lnz��K���:��<v���u����l�;0�Z�(�5�~��]V7R��ˁ�y�J��]xLy��W�X�+{1��E�ݭ�h��F췒��2���w^�V\J����4��SL0��x�!�>-�bؖܲB6�����7t/`���$�r)�g��d7�|M�I.��p�~[��z�o �+���.́tgL�bk��Ñ���,X3}�|�Y�!������6FJ ��+��V��H2/����>z�+��N�R����|v�@Q>o��~�m�\�	4C\!�c�F��*���CJ%�s؅�3Z !���W�2��|�0����y}�U���!�[45)'db%W�P����+r(���$�0׃ݞ�WQn�����jR�A���pA5e�=���d����=	iAQ\�T/�\���)2����$�m�ɖ��f�r�O Ϟǫ��'�|��:T��O���������Yel�~������N�FK��Y�-��3�`c� �Q��<eq�c���m��}��{����0)�DX �	��Z#N����?-F���^[��<q���ȱ a%�JK�T������K�uiݿa����>�1b�k ��_�J�#Hx���~<X$����nGV�啋�?`