XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����(������w\����%��arE��Y�^�_q�ߋL�49z� [��מ.GjQj̣�Y��a:��`��n��־��l�L�������W��h��A�*Ή��FZ�I��2�b�	�	r.S�V��t��]
:�Kf��_&h���<�L}`��E�◢iv��u��&���:x��ryL���݂vr�Pk����l���)W��,���b߀���g�i!6�����T.��8�u� 6���̃W|��b���T).��}h�g��^�)��� �虎t?��,�m�Tc��ٞ"�~6��9�{M�M��K���ȗ:/O���7��%w:lQ������O� Jn/��=\z������)�4me_�P;�wy���G�Ӻ[FuiFֺ"�[�FQ������(�O��v����ٟ႗�t�g��IGyO�&<���V
W_"y$baB����(c:�.�0���?ڏ�w�]�Y/8w���cE�d�\�F�?-�\�ʬ��o���/�HR'=�P�FH~��/�Tn��|���mlh4|&w��k;�&>#;��� �I�~Sի�}_x��Yӣ��-��.E�q٢��x�L���Kܲ�H��# �c!��% �cGN�P���Y�.g-��"P�� o�T�P/lX/>4 F�	tk�5l����kx����
� ��TQ?�,��2�I���0~�J�%�	�z��V�:���n�7,{��1�I��c�+|В����`��XlxVHYEB    fa00    25201�ԓ�����x��;�+����!�Jxp�=�w!����:��婜u��jrA$�kk>L��]oV�PVPQӻ���h[�FF&�Ѻ?w}��.RC�N�@���^LRNY�����m�$G٣h�ʴ�?��������t�31<,�&�1`�_�/T�Q�	[�y��
=R-z�4]L�-rGe��i��ܱV�ق�*�k��s#d��!:�}n�4��b��o۶���JW������'��=���!dC}��KGc51�
�8��p#��� X2y����6w���][�6 U=P0��Z��wp��]E�#{\
o�#����T��gM+��WK�9��1�@�qq�Zaն}���NP�����0�~�-M�
�/ˏ/�|Qq^��BD��5���\�o-h̗�U�/���14�R8�"�3������x�[5u~��X�Ȁ ���<����k��{@4�ε��X�`Zs6EiH��.pN��ԯ�̈��½$�z�^V�h��yf�Ф3.�SN��K\�8��>�]+�"�U�j�f�Y&Vh��n0 ���;��݊�-������)���';[��aGI�E�c�޿Q�eN�f���4z���1�4}�f\'d��'�(���������v�Ml2�V�
��L�-p�kd�ɐҵ��i�s��@蝇�����2#��:p(��[vv�U�F��+�%��IL����+ �i�������^DBL�s��%WͶ�Z^��q{��U3���Z�6gPUx�ih�| [�q�Pc�glX�8�-}ΐv�p�:�&E{�
�C�A��;2;��\WZ�N���rKC��z���)�X�G��ђ��1��|�٥XQv`{>��>(�W4<CX�s�ش���8�j
����F�g�Rh��xY��ND7��	�ّʧ�*/�j�r�4�\8�6\�Le�%R^��Ž�Y9�N ��~����/����1)�[Q&�mW�5�ܪ=�}� ��	�9������Zmy��rZ�N�X��0��2dor�6L�xXm<�o��h��������Xԭ{��&g������ kٵ�\o�W�hZ�ƁDa�b#�E��������o�UY��w���,�p{���MF>Z�|�uyOg&?"���>�3�-��g�/6n�M3Ogi�n�rf�O2)��0�3*����<�y�6 �f�BA�Z4%�_Be<�Ǖur#�=��H���|hk�'�i�n�Jm��S^U��K`�	O�4Xh�h�>U�0
t���G�i�&F���W�|O;ц^�cI0�L_X��%��Va���7ml�����9���L7�;����<n��u#�z��呡�8؝��i�N���s��Ȧhe��ψ�a |�@%�����a�-�)q�З���Cζ<�6()�?�_�#Ŷ����T�+���4�/�D�U�رQ�Q�Ҭ�ϳ�׼�;"?�0jH��٫��J~�(Ų�؈�1��g�U ;h�fz�~iZ��/�Np 5�}�� ���*�Z&�dg�����ژU|�enp��Yk@��,�!o)PB|���e�6��s-����q؁���f-ˡV7����,(��徑�?����煅)II{�}wp�����Y�n��U�����^d�|���S�b?E�y4T0Yu�J��G.�N41�"���3g�<]��z8�#�Hӽ���?4(j�.�y9�O8]�)��^�D�B��� /��Pw�9���j�ѷ�܅�F�]���da �����)<^�֯�;~�������Ɲ�2J��đJ-��<��Q0 )�z\�_�C����,�;)�H�8���}w�T�e��uf�NoǷ�6�"9�9��ȸ���9�ћ>X+oBD��֗�	>]��2��3�m�C!%��"ɲ|e^@lfܲ�C��1� �~��o����Z��������/��T�ď�Wʙ26��7w��> ���OƠܳ\�g�b�-������f2gc��+9����mZ�V�:�D�z~	��O8�g �h�a��q1��J����F9����u���D-y�$�ǡ���u�� aB����T��Z*�qqdr���R1�E�	񱸯G{A��0��a]Q[Fg��{�ܨG��Y��@k���6� &�J	bX��z��d>3rC�)?a��HZP�����C������ ���${v������;�>�z���P� �aw�~�@V�ܖr=i^�^�NQ�zk����z�S4�gAǍ�0�:6wp�nc�{ݟxw��P��#C���:-\�z����^�Z���P����w�
���\��Y�gx�K�7�,�4���T�+z���S���u�+ƉmѺ�uՄ�Eh�ObI1F����"���h�a�	�������tr��Aܔ�`�1�@Y�*\{�cr��a�7q���VL�c
�l���q/�DgČ���n������,��3�f�9]������B׳�<�a�7-�%a���q!\!��#��*`0/�o0�T�u
�q 1T���Mθ-}�%�)�9h�;�(w|BP3�/��1u4u��H��w���a*�����냮����v��1B�7!#�O�};����-��=��7�^�R��$�6�7�GRo�<!-i���;���<O���R�䒍_���҉��W�z�Hp�"~�p2�2u%Z�Ť��+G ���@x����\ው�[�6Q�Y��Yj������z��I�2�����tff��R=�kqѓkm�r!N`�-8�&3V�@����r��YRӮ�
�˖��ѣ�S'��n{�Ϳ>�����nX�g9�֐	��oGڈ ���{�4�l���|�+)�Ɏ,�c�[p��¦O�
XO]���m?���؊�%��Y�9F�S�@CnqhP:s48坆4	��`�d�Za�ѐ�0�R�ٿrE�]����o�G$��x�;��歗�BU�fQx= �->[H-ˋ��Er}��,��i��-�>EEA����nU�i�Щ%d]RQGn6���1���ԩ�bL7����,zu�wV��y�A�C�=yF�rK�����*ք��C�<G���jPN]��V3=-ƶ7-�v?�qN�H���]$�U�^�8}c����?�<� �8�@0q��a(�e�~dh�_�4����x#�?t���>P�y�U9˽Rv3o��B��'����ҏ=Txt�P��s��}�u/U`Kc<
��ban:���	�hV���1Ě�kHc�t=b�f|��w@��N�2��N}Q?��&����P���4��`v����F�7�pDtT�9��~�>�q��:� ��M�'�.���D�������9���s{4�f<G6�?���R z6"��'�^�1�?*��{�������{ߨq���?�,k�j� ���c����1I0�) H��.�ϯ��� /���M���	^�ਰ���&� 'JUS�R�,b�
l��s�͙�I�2�8#��֩,3]D�z�(�t�-]j����>�u;
�p�*0�awW�l�*����-oP�"��D3;�Ŝ1�J��I�6=T�C�x�ܑ��F����)d�-*M��f��iӬ� |s��#��+�ŷTg.�9ʤ��6�9.L`2��ET�^a�j�I��U����Sl�;8:������9�:L���@)��xu��'I��&�!�Kz���|��wP��L-�q�fKuce�~{��׼)�]�!b1�R�B�͚:�x�dI���ZXm,��0�}�����&�9ٌ �~�%Eܙ���I�9p�ܪ�?R�q�VQR����Ul���'�,e" {�����������e�^
���D��w:$E��o��>k���k�m�	��g�j`��xE�-	������*���^ϣ_��Q	�^��"�0���z���l�_�����Q�'����;a��2�<r��Ȕ93�l��D��31�G�d�Q͊1Pb�	g[t<��%��r�D�J��ٚ�](�V��3Ӷ<,^)�����E�K�o��|�:���O��s]�h �h�����t�Ag�u�38���nH;���a+N�N�9���]�<Df�ܶ�����!�X�4�)m��l����O�d��?��\C=���K7���7���t�/�#���;����L: ���5�����X��"�g� L�\��K�?L<�jP���CwЃ&�]������C�Q)��}vĻ����"��%n�%�7(��X�*�|4x���sc�O(�`����1�?�<��q���q@{y�B�)�R���6`!�Bf �6��HUo��?u��V�}��"��^ܛ#U>V�ܐk�Ls�	�D�cD�M��
���"��<�~Ifr������/c?Si	=���ܿ+��D7V�*㰒� ��YTa�U*0fv�����_yG����w���٠��c��_�R:�����|�]�Q�R���R�gu���sfZ�Fm���u��R�M����qySy�iF�\�ԏ
�=����*6�n�é�v�d���[�/�P2<�I��jf���t���H��RE�!/D�G��mb#%��(\�BC=
qW����}���������e/O�D���R�U�2{�S
��!���)���c8��u�� �9l �p�M��$yi(Y�h����KYt)U�z�]B���_��p�cpXAP9Q'
X��]S���[�{�۩�5p��ٞ�6T�F��o����n� g������Iܺ�T�*ٮgh�QRQ���nN�a���}��v�윮v/��U��;��X8�dL��1���&Lp�k���G��[�T�,˚�c��2-i�
�k�=I(��X���jĭ���,,h̹ى���̅�ڏ��:�;�}~��:�h�T~��k�)a�����0���	C��՜g�Dpgj' ����;�<���!��B�ò�"��jI�uj@,�jq���jjEb�5�*�X� �^%��'k����\51����uf��4�6 nդ1 ��]���û���c����b��=�����cYV��J�r����)HF�R9d��x��#4���$]غD���B�y��R{6��i�_�7M�Ԍ�z��֗܌��u!�2���fq��*�ݜ�t�(�i����
f�x̵��K+f�����ڠ(��G�q����#-��� E�ݺ�O�M�~i6�>5UY�qծ�s��& ��Ӯ8}�
�uf����1�B�a
�wYc��"�|M.�$13>ˣ#[ R�cr/��lP�`[�9٠����6�It,:����/��#������*�~�ĵ�~���4&�d�=�Z&Y��� �_�:I�� ���#�H�ɚO7q{įM����m�s�]�k�\Hz�w�^��Х�(��!ܤ���UV�E���X�7y,�~WM��/�����p���'������^�[�i^qS�X?�z�w]ҩ �|����5��"C�Q�7 �)�%/Q��tr'��2	�� *%�uT�99^I8��_($�R�Y���D�x񧓖W�U;�ڜ��n%�L�EB�©-N|����B!�=�F�S�CT�ҿs��4%ݞ�T5sk4w	MS��nEк�u���_�T~�U+,4��QjW�-m�>/[e��o�7�8�kʻ�񇍥�2Sk�/���#�K������W�-\6��'r^/������My��<c4��SU�(Pp��Z�\��[ *��� R}���%h��a��r��)�����!'���Bz������A�'�?Z�#�-B
�$�
�b����?l9D��+����A^�� �Z��/���������a_����!�$/[�.k�`�u�D����<�
��2�}�u��0�aw~�*�M���l37<!zN�#����_EtHڈ��$�c��7���ki��ת��<|<	6-0�����J�){F��+j�4�V���4��g}�*\
�x���lu�Q/"��F�T��m,�n��c�F9�x��	�N �ʢ��)U���%8hMO��#��y���&0ɇ!f��?/��)ܣ�@�����FƢxm�y��S=���HX�������<�^������8L厯��P, )����F�e�����z|���a�*T-�:['3�y4LSᰍ��ӊ;P���7�M|m�I�[3��9/���4Ǖ�G�.�� L��s6�lN�d���Q?܏Ϣ$�~��f(����%�U!:��b��c!V�ԛ�]Ô�	�Mt;���Z�_�Ko>;諸{QuԞoO��Y�L*t]��g��v_�����L�*�/V��q��8�$��	�������w��g*MI�P�@��.��(\db�bt�hy�_�z��dV=���k��lDYA@�:עQ�Ss�4T T	�Hx�V����$%J�|���S���l�ml�ߑ�]0��=)�O9E�m�:��H#̯�����9Nu�b4/��D�:�"ƽ16lÑJe�(�p���������㈸y`�,r�ߕ6b�����Ko\�R�_@3�n�a��Y<�4V{j�;ξ	ܪ�k�6�F��6�V�>�-T���"� �����%1�YJ,�k@�*}"�J�б��j�k��%5ʴq� �>]w�;�}�mFSR����@܋���ݲl�}@r�Xm[�r���I����f����%^y�M3�v�k����N}�@;����G�|������^��|��բ�O������>�@@�����t��cn�c��@�asZ3F�r��v�]ɟ@E�R��SJd�eX����QG_	S8m=/h��{��Hk�kP�*�������c'��شG0M���ܙ2��/(g�|4ˋ"�S�bU�g�}���"���8�!�fUQ�7$��&���x~������t/�Ԓ#��<�m���TY�����;�jc���ω\&�_h����o�Hc��_�_����l4����;��/ć��+��?�W:^�����d�vG��r5a�3�3�B�{�����F��T#'�:���VΨ���Tw5��@�I@K���)L�����UtH�\��&����.�]Sϵ���.A�&G��L���9���ը��i������3�?�pFkbz�]�����$�Й�%(�5_���0��|��^���od�y��K(��4A�_Y�٫�^�r�~��<�R���W��,�伆*����d���TY2��!�vO|7��b=���uV�`���v��"w�t���/Ђ�w�t�y��n�u%�� .4�Z4K�YٲmN���5���Qlв����H��:N���9\�B�Ax�.dZ�S�μ��D�R1������N��=qAJQ��M���D(E��g	Ñ��m�i���9\�$d!�m#��t`��d�&^�x��3�Z%�Ǥ��ي|}p�
��jRg��Ur�f V	:dԿ>��=�-�<��!蔬���Ⱦ�}d�Fg��1�Pʪn
�3}<�pT�=c�Q�\Et�����2079�x)������A���[�ѨEa [2Ox4� 6�����vս�_�P.���� ��#4J��ff=���0������5�`�b��m����oqkҥ|��C��R�*$T5��p �)�.L���$�˷��5R3ݺ��)��~;����0��u�^�<8�v���9mʽ�אf,߬�Y��s��0x���aƫ*��CQ\���\�6FL[�����<z��C+��Z�,7����Vf9����+�-gN��k��x�^|(�*�Y��I���6X �0�(�#��V@�*㉋*�^���:Tr�=v��fqr�`�!���خ-�`���.��%��N8�6<�K�����U�E���v��lH��گ�s���ڴ�6jKsse���rq,�����Ĩ��>�{�a[}8bS�O1�
�@��{�KGoa�2����m���Ԃ\+v�z�9Z��W��j�2�P�;z��=T�wz�l�ˊ�
�2 �%m;�C!4b7�:+c���?���C�ˋӗ��Q	���y��&�=���2ޥ>9���ZnyH���q�YPa:|�ȥV��f)�V�0C�on?=�#�����=�+�OR7����y�~;M������cT�I�G+�&�`�a�|]�\�P�ٔ�}i6����h��A�^[($κ����kP�f���6P�:VƎj�#��3�T�o��Mm-�#���6�5�W[0�c�R_�����ӏF�a$�5���k�١UA��A���;h�՟C��Ibf��+�d��\V���S��#��_����z��r̿8�г`���1ꜿ3��S��fr��=쇈f�u[���Z�4[=y�5+��o�г?��H�����孫e����=�<xr�Zo@S�������o<>��g��>/+�Y�ƅ���u*l����@��`b�����#�����^s���~�3�6�N_������ zX�k	��4�/�g��Q/�=��wȥ�HG��i����r�o��eF���N����/f����fX��~6����U�����y&�냨�E韈��e��I�k�2*&1��-��Hp8h4���n�w�ql���1Ih8e܀8/he���� �ƥ4	(r�!)}���#�-�������@W�)j�a����o Ohs�i~˰/�EF��*_6]:\�IX��n�|��7�-:�r>
�-[�q�'���2�}/(��}j�m��^�@��������,NY���?PE��!�p��8k7���.�K�t$��(�	�&�X!���C����j�P��@w㈷�̴��~�`TFK+G�?y�h��{�d��-p����K#
�
i1\��Ѳ��*a�LlUdڕ7e�ľ�[܅m��~�8²��&Oiue�4�t�f\zJN��7 Ibo�_C<L�����X0ՊC��ks%��eZ���r-���`m@�> M���2�+�b�i�s��'�iT'�*��$�g~���b��LQ��펎6y	t���a�o�{q��8$�l�.`��B=j�7	���Ũ��5�l����0;�>���D�Hƍo��]m%�\x�)_�3k�������2{h�q����v4g�,)�Ί7����Y�بɨ<ҷ�ǚ���H��)����s����9]RU)�c���Ѕ)�M�����݌�!��ܸr��g]8@��G��֜�U�L����}5���M��v$��t�z�Q�a���ߪ�d��bS���vc��A���~������wڿS��16E�C6�Oxz��܃���4[2�G�9��տu6�����X;���/\L��r��1�Q8��07�&�bt��τ��m#B��`�¼
;T�i!�U�*R-�L:���C�;y�<���T�;G�7�#�ϞXlxVHYEB    fa00    13e0��7<��]��g���i@�Y�Y��K7��c��
��5� @�֌0X�#��s��,8K�����`+|!�y�P�AE���v�d�	T<s��Ց�<��M%�y�Y8��I��p�*b;3Ù'�3 'u�����u(x3	�
3��H2rz� ��G�Җ��[�����g���"�!�-��d����w/KTR��$�������0;�9wi���Q��IiT���Jl�Nt��tr>#,����o���m!g���	�F)�o�P�z�Gd�������R("%k�����9�ޏ
� ��/-��k�T�L֫���=�5>��8�����g[�e���a(���� c�J{}�LoU[��ƶ��
;��s�)�!��
�u���#5�����9�Xtk��f���x�����IO���$����x�{ @.��9��<�rR�wG<[�/��^��:�N���h���qϜ[�Yd0tYCv��ɽ��߅��ZaQ��	网��R@���;v�c}��p�2@����*�'@���k g�I����3ˠ��W�Wo����_x�h\5��3�~Y�����A�2�q�Ά�,>��8�2����V��D�>�?Ԁ�I�S顶�QS�8ny�CC`+!$�3�M�Y��2��$z��8n"�[��@�Kf��*��=.�5i�¼Ί��v"�h�B�h]�0�PT���f�,m$z�MH)�Q�Q4Č�D@����.
��+
M��(����l$�9%Hig�����l�x�l%�r��j�j�_�C�7y��*e��+�A\iP�sT�伏A��YU
�R?=S�rĐ��3v��c�j���[;��?3��BԾ/2�7�0���t�#�7~\94ės~p�-��e������Sikk����*�U�>ޝw��������� �~Sk�]I�i�=h�2~/MZG����j�%�-�z7EM�c����,N����v	ȱ!�US}pd8.�@y�����J�Xa>T[�h�3ա5�S�a���{�˒��4����3o��	� x8���|1��Ń��Ӡ_s��߅�G�P�:R��	�a� ���#3���8Z(�u�sV�dq��/3"]���8"�����/�g�|ϛ	��P�0�$�9O}�p�ی#|��W	�:�Zkr&,~��JE��x�],���_ �F�a��@�L@�QAX�~�]{�w��<\��ݠ�'�B-����1��=�$fJ��@%�5�
�BI�'�~@�l���+�ly�w����[�}㰈B>'�x^��h���L�Dq����G�$1y3��v8�M�CE\wQ�$;�%�)��;�r�F�'E��A�8V��v�w��7��I�k�� ���h=�&�KB�G�zR�o9��_%�^l�\V!Z�c�&��=��F���'��+a-M��f��-�~5���Ϗ�Rԝ��q6x&��DjLl*c`|qa?��{>uw�`�Dd�b�3��)�����0�d�nN_��q�9ЂqzeO=� �	�Z�{,BSh��>��)���zpkGs���#�c�z�a*>��ū��K9a�ܢ���ˁ�� �9�v�}9��V��;��P�r�Ƥ%�[��,T�N�VT@�XsON�ê�ɑ��Q�����\@P=��V6���2�*޻���r��d�sX)7J%=�����M��Z���>��'*��Y���{+���S{twm\iA���Nco3[�J��G$ն|.f���)�|��Ӳ�2%���T\��q�D�)�B�i���8<���w/��(��!+L��PA�{Y��0>.����A���t�ZX�Bi+q�6�3dMǶ��9WU@L���m�z���rdk(�r4L�MS_� �!o-��DF>?�u��G�U�V��9��hym����k�)c2��t�&��C`S�G0cCrJ��ە�C�:��7W��������	���/�uէ��?b�o�5�΍�I˄��;��d���Xf��J����h���v��`��ǰ��&[�u�Tt��Us�oycxɑ�?풙=��H�>8?��d}7�@*�H�84������U<��OML�Q'*�n�/O����M�Ē�̲wrMq ���|�_H�H$��7��]��R3�-$p.�,���V�K��}��»���o!�azw�([���PF<���@��,�F(��3��ov@��U��i����R�4�[E�$_$/�Ϡ&3��0z~��Y4����a��]j�ځ;k�42U�`wbƎ	��'ʅ��>"S7��FH1&�n\��1�6d��O _���6A$���yݵ�O��e�\t�^?���9����@qD\��^r���nG����O�C��	����̈́a�!wC܏���l?�r"*G�}���g�e?,/AW��Ν��Z)�6Qy�/����O�-$�7��If�`*��y�<��i���
O�ތ /��}���gp��.A�O�S�����s�HW�7�,�U*H,�=M[/At�Z�ձ�-�=����^���H
6Gj�-�8��+�����5%�RX��ͥ��9���R�R����b_��^�����7h\���š4���W�,nxN-�X�q�Q�p�:0�-�8]��R<�d�泌5���@��{ҫ��l�4іN�ـ�8�
�E�	h�r�/�~/�!L&y��?%�����1Fd0AY�f�Y�~�gL��=����� X|�fS���;��1 �p��a�0iڔ�ڔ�*E�vߌ!��a��x�v &��ǣ��x���Tr�R��p����>0r�)-��X��A#����]'w(�<~�Tͪ�X�D$csU�֯&�٠"�R��ȵ��l&*��-�ૹ����U#�5��|�ҍ�f�Ş|V���L#i�%�`J�Z�	-u��f���*��ćA@0H �G�A��?��8$���p��-�z��l����*9m��J�`O�`��F?��
��Q�Վ�����S��,re���h���{����_�EW�r��� �zh�z]E�����zk�ER�e�&�4s4��:^��-n�ޞ^6}3P�tۮ_�K8��P|�a �P��Q�������mU�0�ᄬ޹�^Oؠ�2TO��[�?JH�ٍ�`��u	�5�աѡ���e�J	raU�����ǵ��r���E��PJ,2�J�L$��GC;���7�Ӱz���P*��kJh3�F#_M�i��W�6��qO�m���Wm�5l9�/ �4���b�,B���6*��e�r�i͟��:I�4�8?4<7���}c��V
��&')E�w�.�ԝ���3n�<�l�2Q�_����g��5�}b�N�q��#�����o���W�|�h��?�-�-�i���6�Ӓ���Y>�66�i���C�5Nx�	�c����/l��lZ��p��B��`XF�����r��H�Z���j��hKU�D��s�a
H�/Q#X}�j7�%,0�	�j*��p�OÅ�{-�M����gx,]iԊ������|m��0�:�t�xjIB������_Ⱦ�`h��[@]F����ڸoj��Q�3��qMT��:��	�S��s�˾�O��J\�����8��l�G��Sۦ���;����G�Ʃ�?�S	�xLK��F]��,a���v�X�~I7�m����cT8�����AJ�A{��*��"6��V֜�rS�N��	�¡��1�R��;����~ ���W5�qE��i��r%���=o�"�Ţ���̚q������c��[%Zh�"ⱔ�$2�[Ꮒ8� ߟ�RNh��:�괇�����)��F�c�jD����s�l�p&\�5\Ԏ�ؒGl2٧��6�*�����)�؁���8��|�������< F���>�\��XM=w����-���d����2�H�7^+1��e��֜���Lg�l�62}��Ȭz��F[���W/�0�I�פ;�Y��7��n��p���`i��D4C����'#M<�8�D�D�@�L�gA@`�	�dz�P��
�T��)�s����zQ|C�3e:�w˛M�������K�/�61��O���Cisi�9�kn��V4Q�1[�8��xa�Ӊtտ"�����*������`�~A�V��.�y��6�0���Op@8���T�w�x��g��M}U�� {��bm��砣av�ë��殖�{s9�ZȭTy�3pˆ|/�)<��7֑(<_�Ζ�� I:?t��/�ǅcUI�[\�w#�_��,EU��f�⥔��v�!��-d%�6�,�hO$}L��b�W��Mħ`;�놕
(i�g�ߪ��K�M�A6^mJV.{��P-CIs4���Аa���)A�=RQ2�
;m�h�G.K����%O���d	��R�l*�m�����b���2w��N���\\x-_�*��A2��b��+C��p�S̗ő��Pg(s���l`��^A�;���I��$���G�p���p+t9�����@�
-�_�����dY�j��e߯��j����b�p.�/3O�8��2P˗�k]:bO+Ý(/Xz��������Ο�7Et���ͦ�Jn�x��5\��⏎P��<G�[�d*�$wI3�
?N��PEf5'���L?�\o�aӲ[����/�J�x��;D��E�3�F{7�*�7�A����
�*�r�D9��S��jki��s�F�-]�����
�9%�*�
w���޸zMq!�u��Z�E��������S�TVr��W��yl�S��gc�!�K��X�� �;B�v�l��<ۀ��FR��[M2������C���b4&>�����D] ػ��2p!CU�c���|�A�}��>x��Û�w�\\����u;�Q�o4�%�ʃOx��{�uK�hJm,�Y0�w/)�z(��0�4�E��)뇈����DLf���^�5��ꮳbȖ���ޮ߀�<�3_�h)�~}6uQ,�|T�<�(&y��
P)0����3��T���h� 7�#{�� 3���p*�������ą�H}��$d�j(:�p*.�@���]�XlxVHYEB    fa00    1780��m�??3�ڮ��</�����y��>��f��y��$�g~ ���鰎���ᐈeN�2�g?8MC�,��Dǩ�j�%(<�/lR�Waz���W�d�`��Ĳ�N@�k����dG����@�\:�%Y�T�+mAY���Nm��F�y�l�.
�����q8�O��|w��"d��%�����y&Y�&��q�>�)�u�;l2�>��tY��3Y�C���N�me��[Uo���PB�+S?�@��R�v<�*+_�q�f`2 �Q1��yj{Y��w���3zv�7���"�/O��?����#>�w�C1��\e%�=C��Ζ��.4�)#j��Y!$�yG=�܃<w�vE��ڢU�.�y�����V�h9��Khf���t��-�lXuw�\��0T�ת��k	��E:�#I��F��zǅz�?iT�sZ^������H�s�YQ���PܷS<C7ū��.jƧ�c#�d��������H��Z�c�S�t�:iį"Ш�9�y�P�>+^����T�ņ]��>�ݬ�*�I�� ���PlY���ę���0̊x3��#YL+�x�'~�D�u��\.���b�C���]��5зG���E�_��9p5�w�dr��Y��t��#Z7�h�̍:�ʈf���m���	��z&��a���Qa9]�~�)�����zgY<��������0��0�˒����"�;c�����;j�ۼ��]͏�ԉ\Z���\?4F~�p�b=BH�E��p(f]fv�U�f�<4k`�]I�p%C
Np�܊i]	,n79�G�9�/f�?d���M�M�H|�¸j��lF_��	��V�1���K�o���eN�V8/�'�^�>�w+'+´B���+����/���������T��g�>�������5ϔh���j�-7/hTؓ>w�p������~_�Ҍ}<Z����B�<��^§jZLS_�isb�1,U�vj�$��;��º��Y!��	Ƣ���_&/�M�W��&3��[�C�w�Ǌ��-�����Y���A@�+ռ��CZ~�a�{�'��O;�ǥ3�o$�+�cK��½��Y���"drWA��sϘ����骪Xb�A	����BwQ���ֵs�O�4�q���0jY+J�~:	��u�����r���B��n�h��Ȫ9y�����uj����kNE�tCE!���iqv����0MD�5�g˄:u���3��
t:$�S^6Tak}��Ҿka��P�9�c��y ��'.L'����~ݥ;"s��.�>Q1�h��Mf�	&�ƅ)��^n�T�lr�bhe�~m'wߕ|��i��������qTid�]R���M!z����Wc�
|�n��r�M	e���H�]C M�N'�Et�(B�(�jR����p��蛪C�rK.9ʱJ�G��n�N�}�>��������V�s�>�C5��
p<�&^.H�<7�{�%����ek��´����,e�A�B����7k�O+�c!�˻a�m���N��Fd�ѹm�?��k�� �����ǈ�0�>;D(�1׸�ژZ��j����]��u���V�뷤��#j�����L�����F�lM�fJ���m�����*!�e��G��<�s� ע:?��3,��o]mn�?���"���T��[��=��n����E��5�Υ�3
v,��g�.u��)˺G19x�蔜�ԓN���QJC���O�q�8�A	������j�`�;�a o=\����4�كY���8<�g�2����?�6���hlb���������C���q���<��4�����́5��1���{Q�J�ҷ�@�2�0��>���n>���k
�_��o�/��w�FCk�	��\�N�.,���'v��kud��Qy����N2H�b�L
1s	)�����o��i�)�J74��������B���,B�N���t�*���wM��YkZ
�&ה=1ao(�C���}X'L�ࠝ����S�wFlG��HA�lJI��oƢ��FA81��A7�0�3����x��K�y�l��H򎎘�X���tFU<��8<���RTw��d�x��4>f���8��b����p�<ٺ�+ܢ��kOA.Qa��{c����Q�o�B]��B����lVZ>ӘA��`sø�S����aKܷ�:L
�C.R��Tթ����
�97�'=}�|g_IAo^��_�}�E����/;*��k�:�Z*v@�A�$e9quF@C*�Ŧn��PS�KW`A*�'�ӵ`7Tj�$�u&��x����3�7~hg����$�Wd�6�((�PF�8CS*�I>NV,�}�����`�h��_hSf_�dFy:*0D#bw�}8=�e���y�<^��PX�p����Zڅ���7Ve�ۮl�����u�����r���i�x6B6+��S`֌{�J�f��� �Lv������n�u.!��x[��V���m��uѰJ�A<}�m���q������J"&Wl�g��9����(�����{�rEԄ��>����گ*��&j��#Ykݖ>�(���#?M�?P`Dȹ}��zcp@+��j�^���=�k#��\�is�9Nh���"YH-||���hS��گ��hMP:��!2��Z�!�rlj��k�!.*�x����ls�\��K���rLY]�v��Ls�4KZRlL,�7``�����=�<��ǈ�
yWt��[_�~��K���d©Xz
D�z��̧��k����<k�6��V�V���Qx�ƣ���v�m��=A��Ndn~K���wV�C\k�dɞ�|��[T�.Uj�AQ�/Xd#�)۷����!.�sӨ3p'v��������|���*'y� �B{-lV���!&�՚͂�@@�x�m�\��w辊��-� �_�:�l=�117]=�Z�OaƸu�W�3�%o����+Nˋjޚ�H�"!�c9��N��]��[�iw
����^�Y�f��
˾>��nn���<���-zQpX8�Q-��T�I��:zNΐ��R68(:pP�=c�!�O1B�Y�	M~w{����%������Od�
�w�x�S�H��'5҆^C⤜��v����������#l�j����&7!GM�^*&���j��k��"���b^Ҙ�ɛ�� �/�K�Q.`k��a��W�\"�,<$��M�Ȫ�s��ٿ��J w���m���J�bQ�_/>����սd?����{�L�Yw�}j���f�~�W~P�mV�Q��A�����L�SW�M+|����ࢃ���kDnIS~�Q���`��O��)ߧx��Fj��2xiozg~TU�ݻ�!�
��)�d���Q�,���ۢ+J�0R�P�-N�_Ă��O$jEY�G�>}��i3F>T���H0�-�bA�o��j��d0��:�Ζ��0h�|.@s�"��O\��+Y��5�]��0Q��OlB	�x�b��(�жKt#k˧��Tp��*�$��ec4�V �>F�i$����z,΂�!�|�	ƴPA��lM�K�T��P�L��A��򶭓v�fze{>C�&�O�ib��j����9���~�y�dZc+�z=�u�l1ղa�ɝ�I�u�̶O�}����CHl�hk�l�>������ew�"����勺�F�Da@�s2U�Ḅ4���W��{�����<H�ZH��;k<�$W	��If΂�G�_ +��(zcD]0S+��G|�ݯË�ŷ�|����q �~�?������t�$q�o]�ƼL����m�b�wR�&2{q�_$�c�/��0���Xw��=~K�l��0��B��|��C�.#���� i$�x}ا
u�cBY@��Vͻ S��ٹ�'��A��7ǰ���;"L����(���$C���C���f�MpN��_'����6�,"���p�'N��/����v�~֛����;Zj�Wk�Tl�s��FL��@ܤ�OR�=�֎g��b�
�1�bp�:3,��q���$��f����~�t2>�v;mY�	Cpذ�
��&�Od�j�\���Z��.8�f�� ������0��z��H�`��Xj��v�W1q+�ەR�1$���֏gHȍ� �P�����ܣ�`0ׯ_��]0<B�[ŋQ�r�uCQD�3�3B)rHH*�����3���
ny��&O� �X}��FE0�X�lE��"�xn~�Vr��ʵ�]�i�j�7l���+��-.�ANm�t�%�SaZ��jx�Հ�/����$���]�Y��LޅG�44Y�	�{�N/o���
��Wr~>���\9՛�����x�����}cj��U$r�T������֓�̴џ��t��(1?���&E�oSt(~�jN!>����okB��-\G5@1��D"l���.���w�Um��[��SzWi?u�e�~����&C��j��Ny:�@���nt��ys5o�y]\�*"3�pKy��s�GB����x9=tI]���)}f�� �v�k����ФY�V��&4l�	�<�<6Pj蠦NFx���ϼ��C4�S���#�C�(�)[.I�h������֖���'�5�kw|�eэ�!k!���78wzaW^	��Q��꡻�uhH�o��!9;�..�)������Ik;�	l��4� �;����	i������ND6C�朄cI7Ni�b�8�3P���J�)�SP�&�>&S�\=�ϗ��V��W�,t�\ɑ��e0��L���C*�t�lt4�쒑$�c)lO�ddMy0�im0��#@��
?�H�yw�R�ֈ��K3[=�aFz�����e�֬<�P����-)�.0��i�y�k<l��]/92�[�������Z���T\�	�ѥ���g�Vr!�d�,56O9KB|�{M5�Ug���>Oy�����O��-�eo��@�S��� �[��a4�Pl�#��t����M�\��X--��V�+#�h\G�[��1��K*k����P�eJb1}�1�&Z�w�o�/Q"��ޠXe�=Z`�}?��,6�fz��`���)�3��;u�ڸ��>�L�=*b�UU�:C����[͔'�}�>┒Q@�����}
rX�ZP/H����6׃B
S��is�mw�h.�	�Zto'�.��
�SQe�z�ꖐ,�{�h��j�nL� �2ᴐnn-i�q�0/jJ\*��
�mQ�H�b4?��y
��@��6�ll%��&K�[�0@g�K'��{Hf�J~�B��aQ>}xb*rG H�{?�|R/��0@�_2��/@�&��o��krbБ��ƺ�)�Am[�l��`��0��$�4XTxj���B�/	ƴr���~6��9	���.�O�-4�E�4���y�S*HpGv���SQ�F�q����;����ǰ�'�%��e��ء�FS3(��|� �7���
F;�o���{�HD�:�]��0���� ��n�tW��s���b�)�H��M��sG����M����n�VѤ�x����J!��nl\�l�Y;u�#v�b
���[���ޒ ���D�<,o.&��
ᒁ�J<�R�SPю=T���!ߩ��t�ݻ�bߎ�tښ�X���۾���ӳ�{p���wz�����4�`1�����[d��|?��?עq���VO���!�f��p9É+M�:p�X�w���~]7t�[���s���}��Qd<��ab��4�"<(��Ž&�	����'���rƂ���e1����P�R����/����1�G��VFڽz�Ne<�u�vy�F �#����������	�,[e�-�ʧ�o�G��U��$�߫:����96��Z�>t`����Z������E���'.�}Mra�ge����w����	G�C��]xی4CUyN�=��2�W,�^�]�A��XlxVHYEB    fa00    18a0�Ύ��J���iw`�t5�/�S�$�)e��jq�u]�f"����? <���76�G��2���Eڱ�ٴ�=����	-a쳕�̢R4�N�(��0�(����kᚨ�N�{ܶ��^�Sk�"�cy��Qu(�v5:�}����7�L
|���K�l��:$m/�2�C7��$�w�.<C�t��ݘB��J|UP��e�i��*/V�.��I�BpXKd�]gK���������x(r�>���O	�U��=�#��?���x�$o=���Ě���g2�A~�������l+f��ξǝ%(Ͼ+)]�� �����!��9���"rs��N�g3�����+=�.�=��⽨�� �zj���BNd�a�e�{65��G� :�C�%�~�	g> LʪnTi�44&�'3@��ђ����S�;��Xؖ��� >�c�kP��X��(���f�(�f�9�|b��g�oP]k0ǃ8��;�z{g	~��sU1�Ƭt��ekJ��K�ĉ'�3+F�ȓ<��pY�2p ��l$S�t��L�������3�i:甉����_�"�繁��|�&�I�b2]���|�ƍ9ĕ1搴����Z����c�5g�W"CY#�ku)�"Rȼ��ٸJ���ʋ��W{Jo�^���mo���Qs�f�?
{'>וh*uۡ-U�xY&s�j�ك�'���Y�6�,�I�%*��:��	z�U��vG�ݸ��f��u;c�e��W3�����bB ��0B6�i��E��$��l���Pwv�|9j���Q�8A8�h�?��w�8iQU�|b/{������m�
@N'N��?��RN]V@'v�w��A��K!Y�Q��@��AȺ�M~%�����%Ry�+8��Ş��{�� z���H'#�qT8}>VOz3�S � Pr���8Z����ůr`U�_�������#;~�0E)煏�/e��X���'����E~��g��Fsꟹ�:�-�!Q�*$%��J��}��@?詷�iüR���E3�㐼�����(����w�jo(�����K��X�+�02H��{
k�'�	�ӷ.��˺�ڟ�N�\G�a���,�+I��R�m���5��fz�Ae�i�:zn}�]��˾��L��/��Z�V6�`�m{�q�=�H��u�(�qˬ��������A�x�dT^��1��t+0�F�|��������Ÿ)b�[I����7Y\(Lj��؆yU�뗘O�2�c�Ο�ك��`F�P�E�+P�w�q��qύ�K>���`%]%e�t
�F���|Q�-RB��̉kܘ7$�WЩ�[��ũbm=��֤�y�d�k/�V������t8'��'�����&*�����3�LI���'��0y��"4CM��X�ݴԎ����0�7'QVG&�K����Ǘ�%�s6i�k~.��2���]ZP�PcO-M�j��b�BU+����d�÷��2�BiJ��)j>�c�� �N8�i� $�9�;ݶ�����I���[��H�c6�\G�T�C([��o�"��l���]��(S��㉍�lK��XhQ0�r��17��%��ڊF�u|�
�����
���Ν^������:2����fB��N!-��5��d���g�z[@��,�Y�m�m��W���P�i �--ڑ/!`	=��7w����vt�e����,E��q��
j�֫�Px)�4������zfv�tu[��~���ΜE����]##����6A3��ዺZ�K��\���>C��(q~Ir�J޽	`���R4j_r@��txe��$T1r�s����.Ā��ɑv!~��M���+ޯvr#�My��~}�:��4@c��ҡ�,a�D����3�R�h�3�	̀93J���8��f6����=���ǖ�tH�#��bC)@��[���='Y���d!"����e]�co�QU����"| ��� ���R�ay���.P���[	�M��"Z��D��@���zJ'#���%�@;t�ƙ�)Hvl�]ܐ6�EY'��*9aA�C�u�.ozk!�_�׫ǅQ���|s������3n�|ЙT�o2�K���Oy_��F�� �����/
{�)
WҘ/L���f���[�9(����3Ov淝F�(J�� X�6S=d�ȓ�/܄(�*	��s+:F�:;_�5O�)����;/�\�"��J����(S�������k0m@�97���l
¯�t��P�9ac'ʏ�����EHz�ug��f���i��a� 8��W#�<[rWA�P=J�Y֩��5SՇ����C+kthT�/1�|�]�������:��;�៭kA�+�V��7����[e�*�*��cr���SY�I�i���l��(��2Qv_�{����_�Q�D�����X��g*�]j����8R���-�F*�g㰩��G�R���V��L%����ךD��r�Pî� �W(��H��`���A'B��K+�4�̂N����Ţ�>,gP��k^B�R��ubם�b��5�O7���Y.D��k���
�
���iv��Ax�F�$�gc}E/X�y(����Gz���@6��#�mE�魜�(V^�}�r4�	i@B����Y/����k)���ҽ��v��d��k�^=���f!�}Q"rd�8�\�`#���;K� �����I#�4Nk�	 a��X���v�����ǫOb-�P��S��տ,�8��Um�{�<�� �ū��?�a��I�kR��.9bƳ&���d��];��2 	S��ye��4�7�m 3]�kR����Ȼ퀪G�I�A����¹��l�/��C���e���sĨ��^��7�҃����ӎ#�8�Ц� �����s��aʢ-א�OR��zr{L`��j������gdLJ�GZ΅#Q��ݩθ_5!ih���@�Վ�@"���>��Ft3���c�Dt�QrŅ!�zCV��^?��?�]�x�:���ߨȨ]| YwZr����� �a�4��;�ZUU3ܒ�H8ʓY��NAk��:!�[0��B#��*��/�ΙZ�d�e�+��Դ� �I����I��?1^sU=��pR};�$�!��H��**�Bt�1��cC�oiW�L�CA�|N���n��$��	1j�t�Ʃ�ҪV���dO�_P>�zˣk���x��a�y��J�j�&�ʌ*i6���:�Ǔܸ@x<e�I����Y�>n\����2Sn�a�S�5_�_j$@H��+�!��M��(8[��c?$= ��{g�-�� ,���8RY?�R��@=t�I/öߢ�%X�o�-����u�?�Z�Kse��z"��U���=�Pl�vݸJ�}�Ho+H��,��gt�i������k��� �WB��-e�9,N����(��c濺�p6��FxhV�ghO�i�
�\X��4���a��H.G���T�]}���%��Y ��O�WݍطZs�`�����V���<�%�0��ԮD��*�S���'�x1K?���6X�D*	��<�Z��S�*-
Ή' ���5��걓��*i��ԛ�����q�~['[3Ė� �r:7�h,����ñA<�7pY�����K�xP�������"��т�X����	ǭiv�=42�-$Q-'6��_��r�K�wB��;�!�Z�<Z��ÀC�8�2��'om�X�� AU��>�R�����z��8Qot��U��4��E�Mɖ����[㶓6;�%�A\���s�[1�֒��![^�\Y�/�?
��]�ٚ|������*���n�L7�Д�����=�BY��vRh��(��Z}m#ɶp��_���H�8=c�,p9g�r_l� ��y��J�N�HMз�nR۴��{��fmY.HDX�=�>�?C/F�$��^1��c�u���f��)��y����>\�.V~6�C��n���*&���ieBi��a�U�]tPU]5ұ(.�6?QL�p�Q�^H��$L���3����7�� z�8?���Se��	���SBޠ@)x0��1xn9O@�A2��������:�w�2���A��q�w�.~�C�fX�!�u��NBJ��}�a�+ �7ѫʛl�	-��th���~4�����ghͳ�.*�0�>����V��*��%6��j"_����o�B�R_c��;�������jg�az$�з2�����萯�hm|��ax-OF1��0�H��;Y��c$J�P��$�yc󣀾űx�
DJ@�%�,����P;�(����r>�1�	&1NL��~;VT�5/T
��f܂4"����՗�z;��G�r�L�`?�q�T��ѷ�<$�]���`s��/�ü@l�lB^^�C��|Pm^��:��?aoR��|hN{�h����
o&Ɂ�r��J�ۥ�@Pd���/��t��:ϣֈ6�=	��>[q0�I�G&�JvR��v��9�N�{`f��MG(���1�	�/�5̊
������H��~O��+�g$:@�'{.EG�ߟ��!�S���C9b�(s<�B��j��Y�����ʸ1�6������;��|-H����\��C5��c�����ٝ����Ko�%�C4T5�Eɦ�N�`��-X��͞|R�`/@K8���x>R�Ӌ�c$χ��C}#�,&�6H8K�Uf�A����9���ރ^8+�_�1@[���X����&�bq!AI�˪N	'0����L��/��1��a��'f$�YnN>An@n&!E�!���m�@��_�C�=��#�O�4(����L�gChZ��1Ó}���q�x��a�(�����#~nF}wȾ�{�3q�h�?��I��w��(�bj�������J1<�\�6JYl���@�Ϣ@�<�������xiǨ����Y~
J|��[��&�z�B��|��[!��?lI�d=��nxlm�1�
��Wѭ��	�6�fmW�ב�XO8�F���LN�ǁz�B(��Bz��V�ܘ��2IH?!p�r0@s� ���^�}��Ξv����;�E�B��D�fr/%0�2G*d�L��Nn�����P�FJ��.��" Q˗'��gv.�$���vi�t!x���E����"@���ޝϯ� �H�R�3D�x9��·�!d͹��s��jT9 �[��:���>��ܿɂ���F�)�8��*^�Q�������/���E�O:�'&�6�y[�D���""A���n.T�((A��ft���P� �r^?ͽ��0A~���|AL��Gk�%]����?п�w�v:5��S����q��c���+��_�Et7�H`J�ݗ� �$��0��i��"es-���-M�����t��Hɑƚ�CL�aG�ųONՇ�b��Y�f���D�*��T)(x׃l��������@�2�,�+����W"�s�d�Pk褌�wXⴑ��72w�"�E2@
���T-��>���m�qn�|�S|�T{�CZ\�lz�����S4q��>�-8���O�.�u��`s ^�K�Vm��1�^����QX���Ĭ���v,��6cԑZJ�r.R�5�ȥ�g����$�R�X:I��l�K\f�1!��pᘠ!�ѲQ2��l����VZ���|���;Ȁ���[��2���|[��RV��K
ћ~B������S���&<f��8go���*vC_��Vl���4q�B����{��K#J846����7H�b9��e��ӽ�c�w�{K ���E�i�q4B"z<��;G�Y�>-��(b���T��d�� �:�,m�H�+`���6lquט&J0!f��� ����cNFXT�:!�rӹ5|�����НN����2uG!�n)C��m��<������&���Q{�nÕ~�uO����~�{�����j��)��V�5"����������� �����CΩa5/�X�e~F����~w���JY�
,y%�TG3��k�}������I�Kۼ��9���;j�,�������-b
�;�s!<?щ��[%��'�+��7ۮ{�*��߃9	�!��p.�6�YC��1�9{�_U�?k\�Ҳ'�ۍ:g:�Sme��K���vMsSS�;�?�\�<�c�x�%��&q�9@F��̼�v�DK��9��  c�l���]��	Q�¯�.p3� M�h��Έ�Y;�}�O��J�[g�GG�\��
�5j�@��8�1��H�Md�/浚)�_���@���N��g�Y��Y<�'L+�Ԅ����c� N6�4XlxVHYEB    fa00    1200���|F	|-Bz0��j��@W�pw�v���7�,Z�7�րw8!�w�oT��T�o����� ) a"i�zw��i������5��Z�ݸ<�TG=�Ruʜ��F�7�g�r�>��������������[{���!�G��7�7��-ց�@p���b;߈g�S�+&�F�]�O쭓��쮐����
�_mƪ2\�QXB�:�5ͬ�9�uy��:�J"�a����H������H;+Ps,����GŲ�;f��Z@^� �L�/��1�`�����%�$Die����jQ�"r�mD��&nᏮ-[[�g.��O=�u���z��}�ކB}U�qG�)Zw��0D�Ra�3yӄ���4O�4�C�����5@���OU_��D�脗/�{w��P`k�8��k��;���5�1�15#��V��/�49��R!��3�)ҶMCy>� ��� T~B,��9�?m��U��h�2)&i�-B�p��<�#nY_�!H�I��n�[.<���xt��a�I��������?��5�i�=G��4ۀ�l�%&��\�����Z��G�졾K�Ƣ��}Sr�/�*Í;�S�l�id�}(`$�IG�ɘ�n��Hؤ�/�EN��1�']<�Z�n�{f�a�[�{(_6Ҽ��Yħd��h��F�C}��5;��g���2�N�󒮃��K��F����fy鱗�FY{!0?)�#����N��y�P�J����E�E��$&�w������<p�y�i��C��u �����(�h�\��T��b�\���?�y���]W	�(s!+�Q�NRF�L������a�����,�W)��H�v��Ax]7Db	;[��`��ؐw%5���ݤY5+1:�c������>�uX�G�?�.�r�S\Iq{�=MI����^�C,"R�U�Y����G�ep��X+-��PBj+�uut�e�x�)?If��Eb������?�k�Z���c#i ~Х�`�0O�k��S��aQ�z�J����ّȭ�ħ!�_@�8�q�'���_ClT�>p� ��5�#���x�d�a�:�ZS��@��4�bL���=s���f��p��=?w���i�3��0əJV�(\ ��1DN�Ʊ�����o��4���Т�Σ0�Kخ�`_d���R85Zʇ�a��NORptҭ�q_'�k���-���"D�bI_M��j\��_P��� R��&�Ba�A�\L4�Re�S�Ձ���\Ei�ͽ{�7�W�N� �{:�?cŊ���jӅ�`Z�&����}YR�R[jŘ[�Ҝ���e��i��e�������1U,�(�Q`�3��:�R�12PB�@	Y��
Zd�ۭ5���<�V�,4��ֳ�v�a�rc^�톘s�z�Z�k��z_����W�a},^-{�#}�I���
����VX/�R�ꗻw� R�N�'v�v��B)�mX[^���Lʛ�{�^[������� ?�{|ǂ~w����#OT�^��������_`�E���U��%Uf~G�2qc�cxQ�����%�E���0�4E)�,��PV~��`��%M���^Kn+o��opN ���?���z�^��(�;yGP��J)� Z-��ޮ#@{���E	'q�c[[��u�n1�BK=B(��lц|o�x��b���f�X$)<���aV�z������_<�sL_L}��kJ�X�'b�%ҽt_"��`}7>��N�(���C���FjN0Sp��x]˺���tp��:"�AҢX�;��iΪ��D��g1�d|�͟��_�>�ӝ�][j�V��}{U��\.��� ��F��4����ۄ>O`{N�����t�({C����b�QC�*�������C���#G؉9�����t?���W~,��/��]�jE5*t��>�T�hlJ�Õ�[kd9z��h0g�5� ;y|��)���ֱ�#�H#��AV�wMM<}=�� o@�L3"2�5a���NL�}�ݳ-�!�j�_�]R��߭eK-~}!�)��v�[l�V	��A��(H5C��eBF)�D����9P6�Q�^��NÞ@ {CNj6=�U�����Ĕ�e���נ�I�*|_��__���:~��!�lg�JtW�]�6jb��^v�&��{��{�u���)�����i�5��z���-��\_���z,[V4M.O�Z���w%3l�NJ�Idq�n4�\�o����X�猃	�'2�<»,ʮqg-��B��+�OK�/B"��9Ԫr8����ϙ�4G��I~�< QQ��M7S��ٵɗ����]�9�[��GԖ^B|�P{�2��������o�X5�+]���$�$wvM@(�"�L7t`��\z2j�w���!C%���ԉ7aI��Z���V
>�x8���0��K�l1�&�� p���,B���,S<v�˴7k��Iz<o�=>�2(g��E�vֵ6(--���zڅ����Rib��j&Yr���,��7���8{�g XS����LO����<G�h�J豵RO4�����j�	0�5�+��0�B}&~�c�-��B3Y�ѝ���Q"�F�h�jQ� �_�"\�_(�2�cN�0��diOy���f��\Uu����C"�`�{<��&d+/i���:�X�x��#>���>A�ɥkc�,�D��s�/�>\�s?ֻ�݃��X� s�3V�nLTR��m^�<|�$�v�*"�Y$UY/�O��~/��\�8n���(�g�����Ó�Dt�/�{�8UEV=�8	s��YN�8��ʪ�Haz%'�T4��q��K��ķnd���]�&�s/��x�M���i#���ؤ��L*�b��Oz��4LlK�A�I\%������f]]�����k�J?�w��w4_�Q�(3�	e�Ŀ&��0]���0-�M���������ns�涨Ɗ&���8��Vq�L%�6����0�����]#��Dv�*n&���7�'7
�dFl}�(���������Y�V�\�aH�[oT�Z�U�Ncd�Mt��Gc�n%�zC&?ΐ�I$��þ��K�ʰ�mP���q�l)�M��[i�E/�5��nT��돵���\�!�ج�&����J ,��0#�^��W�h����X�՗��F��QSة����Z�?�>�f����3Y�:�Ϡ��3bWi���Z�.�"
$��K~p����*_�'G�ޗ�q�|�_�J13Aal�U���a>%���*3#��*�qC��;V'5;,����|�;�+�H$eim��P��~�I��D���G`�	�����H^;sX��,IX�jQ��=�Y��B�'=1P]�y֧1�	f���"J�ޒ�@%��:�5]�j�sh :x�� ,j;:i��$��?W��N�L 8p;��ϵ�r͐��$H� ��OVҵ�?�\�bpS^��'�y�HU-�a��ђ��nsV;/�����=y�+���s<3��N�G#z�e;��:�0*�2U�>�T[t��_��8+�}mv��*ف��(�hr.Y��EM�-�ZW[V+����\��|<M�^`��>���j.f�ԭ���v�`h`p��4i�^�$}A5D�W�4Ԅ�1:�n3�P1}K�㖭��\<K�tY����6]]��_�.Ԭ�W����uC+~�Z�T݈(�����B�>Ie�eG�4L$�/��
D��Q̜I�:�����,�yA�e�}���V�Q�A�c�$��e"_�0��������j�6a�U%T�).I�,lG>4/��h ��-e:�yp��]XѼ�Y��V���ɍ�D%�19��o95��2rds����,�ޙ�Cb^ȳ�Z"/Q��a(`�w�f�nYϊbV�]���1������-��E}T.v���H�
H� $G{4ۃ��>�-���j��\0���u����kgI��{�1��B��Gb�G�LP������Z0!ay ���#1��Æ1�_��%�c�/o�y1Xה�!�wu��&�Ԩ5!�Gx~|�`��x<� ��&��~ �a��% H���Uy�^�P�m��n���������V������u[�|ʈ��:6��9��R7l0X��or�~Q;��o)�w�bՎ)h9��eI���c�I�Ҧ�ªgːRet��:~��v9jXy���e����`���tg��'&��Zs���}�w��*Y��40�⨺��o�8+�Ls�b�7#�N�������U}@}/���.�dHqB� E�,�s��Y`��n}Y�1�~R������x����jl���s��^Z��Gt��=��j0����0Y&��1�2U��0MB���Cǉ��W��T���v�~��4֐�
� �_sJ� eG�A;v�P+Li68��pPu��r�I���_'��H��4g�1�6R����<�,�fEzqa.P.^����ǣ�����`g�b��������IP�\۔[��î�π���*�ē�V�$�	�0v^"�3�+�����V^�E_z�#��9$}�ۣ	�(���YJ�Ϻ{;��[�9�pJ�1ܝ��O���Ґ������IeY������d�6ajq�XlxVHYEB    88c9     8f0Zi����gҟGV-�lB�F+���G2���	N�})��"���ז�*���l�����r���)�;Nk@�N!%�>7k���摎;@�{�_
�ۻKCTVtn�r�/BP�Z�e��o�� 0�6������Y��_c�pLP�]:q68��a����W*�u�a�TN���ᅸ?�^� �G����Z�Ǩ$J.�P��a�Q&��
!�$�t�*Vp���d31��/���p��t9Cg`� ήҨ�=W$�����D���^X�xµ��Og/W����� DH^��c�6Վ�-�B1��z�c�m�����j���{���m7q[Ԉ�L�����I�z��?ҫ��Ȼ��^M���gF���<|p��	ؘǍg�;N�;���U��p�/�Ya���:S���\��S"4n9=�xI�B)���\T��ܥ���=?
[�9�Q.��y7��t���,ik@I��-�}�6p~����??`�p?�����65��}������ �%Q���9��1u��t��+�.�=߯���P`~�m�?
aC��W�h��cl{�|�����o�%������sۗ���M�"��7�}Vs?��=qEˇ��ۙ�[j��w�MxsQ
Kp|���-�2�ܢ���ZJ"x*�ӔX� �f���J���P�A��}�����	h�<@��ݍ>e�PC&�G��M
�0��K����o�Y����'�d'��6cJ*�\[YB{�.�W���%39����z�0x�u b�?�"�ai�`
����|v0Řd����B��Io�6.8-_C�Ti�E8@.�!8�S�Fӥ�T���{^ƥ�d&�I�yE#03b@��EH��+m���I[�Rvv��U#�C�B���g�d̵q\�J7%[f�6~1��$4���D�� *.��EH����ܱ�`���gM{q��-�>$�|Z�tW�I��MHU�\�LS$�H��	��%)x ������T�g�":�����#�t�с��;���y��J���~oyH��X�9�F���� �Ru!������i��x����'6\������Eמ C��$�5�J-�l��tV��E�MX�`�9e0�!�rqk��je�"_R �'\c�9N��:$�n��� �^�$,�������=?@=���c�QF  &�/˝�k��Q:]����M�(�1�n`��<x��ظ8m?x~���+�QTǴE�<���-�� _�&�և���lqѿ�+^ׁ��jc�q����G�l�]���׉ mԄ��S��$��T5o:)p��&z#2���I��-�=;��Ѯ�D�ɅV ���0<=���ј���q��
�G�U��m�]نL�fTg/9a�AR�^���j+��~�x�/#���om0�4 pa�
M�1[�uYfLh�n�)�f��t����h~_G�]�A�3���Vo�K1#xP��N����F����b4��j�Fa�FNt�:��ؓ��T��wq����g��>�d�{�%�hv���#�����%{&Ps@#���\J�#�X�v���(��vP垕N4s_�O�b�?E������w܎y��K�B�(敶�eK��0�-,�wȑJuI|S�[���e.�%h�:%�nԑ�1w�;��7�4Q�;%�R=���.ck�#3\O���{+�|�d&�����fܛ��%z` p��x� ;���z��+!D̹늖fX�"�P���&_P���-���B����@���_��(d��F:#�|�San�$َUz>X +�%��ñ.��g+5�,@WM&���[�mzML�R4�����gAq7ۅ���!;�1�rK�{R��7�r
�!V�Ok������@q->�L�NfP$Z߶����om�n��~���N�����^`��w��G�aa�$�h�C:�1h}X��+)�G'-�ձW��	���G�4�zu�d��`9��2����a�`���ԙ�bf�j�"�
�q�Z ���Ý��kG͚Ϝ��EK4���v#k)vE4�:Y�Kc	�w�V��9�mۂ�>.���e^K����:C��PD/Ų��,�C�v\��E��s��/q���ƅ�.�-�عq�c߆*+���W ��*�{������KD�F�eD��֘W��-�G��v<X�𧔒T,���o���dx���=`�����dv�bk���)������*z/^7���/�����b�Yi����0Fe�@;�� �6��