XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��v��!p�`�nN��)�	ܹ	�|�-�_dk�(xp�� �I毁����m�~��1>P8Lɋ�2�x���J��ڦI��7F�;��`��<�^2��6�����p��3m[l�:���]n|V�64���a�����fu��G�܇�:�' QU"�S/'�V�#�:\d��w6���|�P۠��};'̢
;d�	�u��#t��DԹ���<k.���O�T�#י�F���˔v~�#OO�N��Ua��cc����JY�i��6ui���eM(�+w�"�G5[���f-GQ��@p��/b�iy�v<\��:��S
?�/<D�d������4��Bύu7��?ۮ�/���1���g�෶���3��,U���ZL	~:Ҽт<ob��G9zt�%㯤$$Lń�X�����Q�iZB�6({�j
c�RC����L�m��$�����XM�\踲�����*�{���܋�U#��U׈�@8\�f�vV܍�x)�l�R�w�O��U�*���˃�¡<H�����5؁�6;b��u���r�):�J�"~��Bħk�̈�22Z��NC�8az�w�J!���"�48Z��'����+z#��-�O@��99��S�@��!R	���>���	G`[�I8;�Ϲ�Z��4��e3�p'ǐ$~���޴	�QJ��Ht�mL.~������O��?�Ǌ�2J��~�=<D��m�*{�������տt5/- 
�XlxVHYEB    33bd     c90m{\�G��#ܙV�m��1[�*�GR�K�%�?�}�|�' �3��.Vs�~��$r�1q��LNizy���^�?r�z�}Wv��,C*F^	�i��k�K>op������p�:Z*��PT�QhA���`)&vTɞ�@��ZYU$���TI��慆Oꯞ�5}�f��8����q�ˣ��O�}�b���e�$�󳈾o�y$Ŕ��5vt�9�ft6��H�D^+�"i�k��+�2&�Q���<H�J4Uز8�-8M�칈tJ�L��� �]��t;�A�GV���>e[�k�ǽ=���cZ��<��2Hv�[�e��i�W����0�X�Q\X���`��b�qd�.����,~��Ĥ�-aX,�e�M%�m3:J��`�r��o���U��cDf���qy�04�B�n(S����^<2&+�P��b�'X���:��w����{
L�^�/ؚ9[	�����e�vh5�C�+w�2f���y��j#��c����q���J�~���Pι��}T�"��y܋����SP�'*�����K�L������8�
5�D�Ct�t��z6>�?'��KK��(6�g{���A����-y|�[>D��Ÿ����N�z��_|h�mp"�iP����fz��1�rxe��(/��|,?Rq\���\�V�g#r�������E;
�^4�,�����a��l�0�yh_i��?%.�P�5�cV"�4�o�U�fW�|H&�N�τmx����NI.o���b��e��I�o�I����>ˠ�xA�`�����r1b�M�J�vr�/������a�A9��mf�B�U�� �P���>���&�_#��eb�6�!�~��O{�.�\Ť7����'���@7�k�O��B������DQ� m%L_gs�?=Į�ώ��<ؿ�#��J���ED��,��C����Aƨp�]ŴQ�~����Ɋ��Q6�),�'�0d4�f�z�C�|�O��;�ϝV�7td� /$!�]ޅ���44���&l�iB�;�X���&�߉�8���X2e?�rf�{O}���9�Ζ'��i۟h�r]0���п�H�q4kL��(|������N���l����Ӛ�;�/_�TIb�+���?�/����prc��ǣ�@�Xz^>T���L��C��o��u�';M��F�S�8�ߠo���Xҭ�g�t��*g6A�#U���XE7�$��_/�B��&�ߢy[�+�qX���?��J�׊�  4i�r�Cmd��6rR��u8@yLƯ��GFP�jZ�Z`�:w=]�C؞6KjE8I�_�0Ğud� ,�)�(���$tL�qeN��:�\��4G�G����
0ĝB��J�*��FN�9[�Q��~�����b��?_����bx��ZT��O^�z[d���r6pFmq�W�-fͤG��=$9`kF+_���Z`M�7����#`N.dm0�d�#�v�r��l���OvCC�HV�9�[$��)Щ,x�)����@��z���=ΣůU�#	1�k9k!������#/96�I�g�M�%ĭ�d~bo�Ϝ�w�d�̠�Q8A�iʀ�L��?8�1]S� ��B�d��<!���RP
�}�l"~W�vJ����&t6֭H�C�R}�P;0�hڭj�+G�ӳ��i&d��ҲO���Tw2�
�|ԃK��;�
L�k� %��J�u��X�C��X� -Z~M�?��$.85X���M)��V���>��b��|®}�Ȉx�'
u:��_Aܠ���1'�k6�B�ca�T �5�ev�I"TR��b�1<�rpT�{��/�O���?/63�>�W0��5,�0�0j*�b�j/��2�I�4Q��3�e�U�Â��q��"�r��mā4]��΂Jg�wk�u���P���#�����\Sx�� ���j4�fMB�r�!@#<8 ~*��ZY}���CM�,����(m|�ޞ�|6�� ���9��Gr|��U~˻J���ꛐ��:ϓ�4� �h ��q/�e�6��+�Ώ��/��'Ϯ}L߮��-��[�|�~7�yr���LHÚ]\Tl�3� �����K͑ h�S��Y3��Z�nZI�2\�v���{z-u�M�l�}!�^��"����_�����8V㷷�:ʾ�uվx���%~�>5t 02ҽ��.�s�`�A!=��aT����M$y�����SfG)�2-��i=&mi�,�d�Y�̦�� z�͓2�V����Wz���P������ZSӳ�nk����0�5����M�� V��/�_aV�`����:8#����[��v
M�J�]��0��?X(=�N�#-@X��N��\�@!���0yt�m�@A��Ax}v�\�~�]����E V�ͨ�kmW�:x~���
��6�	C�@K���?�����[�6rSg�5tg��%��%�x׼���y/�{j�K8ZK���(��>(^kR��-.�d5�F���\�2`t.Ӷ+J1%�d�w������٠�k�����,���U5J�L��E0��1��[O�/K���� A|ܚ�sy��!򕉃D]f��M��P{VY#��X`痿N���C  b�#�#`Nz<��EQ@�Qյ�=�����u�w ��JE��>K�L
l#,���K/#kH��1@p�s#㞽���ML�=�>u�b�^�����t�A7>cz��'p��j,Bs��+��P-�y:=2�����=���� ��yv�L ��P5y������D�8�'A>�� -
4aׂhĝ�j��%NB����U,h�fM�1��j���.�M@_x��®���KSp~�Ԯt��A�7�b!�t��?���T�����~���0fP��2��H������V�F��Uq�(����Fn h�x��P��+�(��]�����`��p�M�eVϿ��۠9?ñB��"���x5d�#�)��j|�$��tO��J���D,�ٯ���O��͋ȃS���=V�q�Dp��2��|�'���g,_���*�`���3��[z���T4>��v��R�L�\0]��#���b��*���ʈ"��I��g� N��lQtg���J����=�Z�z6x�88�p�ū�.�6��Y�����F܉~'����:C.G