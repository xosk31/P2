XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��R���c�F���u��B"�)Q��,q�@��b 﫞���۶���Hh�C�K���'�|�E�o<�QV�o"�X?�࡭-x[J�S�o�\d%�������g�[=�9��lP�G���r��%HEСʹ����V�	��E����xA�~����xz��[��9��f
�e�C�/U���s�0�i:��FҺgD��ɦ�5=l��c�Q�f}��]"�o���3a���ԉA�d[C���pa�޲�s��m�*EXʹG��)? �1�W�g��|�\���Sۀ�lT��MT��p9OF� ��(�UB�琨r�%�.{Tb:僙G3��Ķ��Z�x� L[���ƿ��&e��2��{��Q���u@;q��17U���K��4IiR���c�dJ��>����R��ގ򇭑:�fI�����z�
��4us5l��O3��X�ز��;[�#tbo47���)jŶ\���kDh�4q�>��`|�:������W��hhad@�_ՠw�6����:wU13�؂S��Ā�{�����#�G��H��f�P}|@T��H4��#UIٜ��Q&@��vf��U��gb��q�`>D
UKh]/��	��Ѧ~���L0$L;J�� �������ǘ����cn����&�Ј�G�cv��}|WF�m>��3RГ�M��E�[^���|	���Ԡ�k�z�Xz
q)���˲P9f����l�ˤ[� �t	�`+�%:�j��7���� �� ի�³XlxVHYEB    17c1     810��ܹ��z.�-�����r�y #��vKB�-��]sQ	=��n����'�]���t�T�	Yܬ���6e�h-lb��7Y�<�\q�XU"m��
1�ӯP,�Ӏ�v
�p��=�觌�0^�|�^m=��9?e�C����*��FP�e]��T�,ơ�6�힫Dy�e�z��Y;��{6ѧ�'!�
��������	���O����������&� �<<=�:��v�����A��"�~�S@]���e�h��p�,��C�2K�1$����@cl�z'H �)#�1H�$U�}�.`�u�2��.w�FA*V�����wfR(�<2���"��L�.�5�è�t��UBچ�>�K��l��*~vٱ�3��t���3��칌�E��ĶڇG+�W��R$�#^�:����U�o��م��ܨ��1�2�DT�k=�����dlX����,C��ɂA�D�2���2_���H����0zWގ�A
����w�F�����Y����m4֚���׳%�$�:Z6��ώ�ۗ��:@r&�|��y�׳���Db�~���(w�S�3��\�R�";'L�y�9��LD��O�������䤑M�h�Y���0�'���FZ~�9��&A����"�m��K�y�$�ꖞ7#w����TA�Ig<�ڊDO��g�7����˒�mE��^G��!�|���e�4�/1�J]�5B��G3��GN_���/p ���)��O�d1�a��a]��͊����Rd���s�+�O��Q+�j�5*��ʣ�D�C����	�6V��S�l�����F�U��l��9� �Y�&�h�t�:��J��qMoy�7w �a��+4^eF��e,��ז_ki"Ѡ%,��	��ϖ?3�ύ�N���mY�Q � �ny*?(�T*%:��O'�򇧵�lE�BC�}�;��@�?{���T�UA�"�
9��,B�9Z�����^�����*�t'����jאg��[�b��|C�Dg��>�F��Z%�kC廞�g�V,[͏m���A֥�+m3v��)XW�8��.���	0b�	��I����=��tܴ�ǩ������IP�K�tw�~����y�O� T��:�"`� (m��*��tӘd���j���={'Z-;��we3K�E��'>�I� ��#��ñ�iMT�_m4��ΐ��C�}�K�+���.���X��,#;�C�|��rb�-�w�0�'�͊d�:kkC��jih��[?V���r��Ƙ�0�C��{��'�f��ӑ@�As+L��}��Drzws@�'��&ho o�)|���/xѪ��Y�M82	3�+� �] .Q�s��sl�����x���3J=��X:�1���i�HF��3��~��ZZ��j�ז���uP���v�}�(Ѧ�{ǖ�FG����ʬΏ�u�Q8g4�C�3��=(���h938���'Dc���U'=�sm�Q��֓ʣ�[�E��.��y��鰭>L��`���}����L��% ��('.�7!��*�zxq�st'm����_�2�X�X�1io+�l�L������|��V��G��G��	7ݍG�A�G�`���8��k�gXS>h� bM7R�m�U�.&߰�)�d�^����G�\�H�\�~Z����ZS��5���|Zr��$�@�rC�U�W����]�gG��� )u�PZ)ˬ���!��������!˓�^�#��L�˖�����bi�����=	l%7Q
�[�C��O��ѯ��[�ʓ�E���+m��	�&HhR5ڇ>��~7Oo��iV�re!!�s�N�<�nV�Q���k��|��w�e<�(�m�b��א���
�^oX3���g���y�?�Zv{�3�a1m�*q���O 	C�³�����k��A����O\��!�)�Cx��S�~ߢ�X
���Im�e0�(�YD��=��wT���D]s��{��t�}�g��O'�<8�7Q>>��,' ���O��J��%�Ѵa~�8���i��2������>���}ne��#�V