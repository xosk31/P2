XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��1�_'�����-����%4���x7�ߓ7U"�#(��H�,��U~(��U��ӛOV%G����o����?�+����w�,X	����e�;�Ś1��:�����D�>A �A8��"�!o�B�����I��ʝwJ��68?�{�D������}��kCqd�e 6_$�}j�F���Q����2�l���r�Щ������Jre��y�6���|�3��k��7$��o=��:�g�]�	�FXV]��O��@���v�*�z�t� T�5�t�0��	�3��aI>c��M,������L�rۅMv�����LG�)7T�����'��p?i|lI�J�H�ƕQf��X�鿑g���eZ3���b��qDm4��EO�D�:Ou��Z��:�4���N:]s�*H�53ܥ)����$�J9ﭮb�³��[1dE�fvPU���'���^���j[I}�0��Pmj��W��\JW]e9G�1�HC+��A����	/�I�CY\�5�H���8q�}B�����{|�lL�;��O�M��y�-ޭZ���Ѡ�8t�*�g��*8���;�y��(Z�*��Q���%(��5 V��T���{ڮt�f�/�҂�w�Ҿ���#4�n��{�R��7A�Љ�����f����/ɯ�p#�§�V���I�����WL����i�pѼ侑c�|���b���#�v6�@S՞��(u�����#�Tk��[��L��yK�7�:b�[.;�}�h�Tl�(����E.�D�w�XlxVHYEB    2cfc     c80�Ϊx����'��{=%�A�菔��P۠�j7�b[=ɕ\S�'��2����f��wY7|��Ca��1/��+�+��}׈�O��
���-����*&:�u|@�(�MC=Qs��s�wg���|�ԓ!:��g�c�`I�|��e�j����w���v�uG���o]��d�;k$�pj��)�!��6��"��;P;,Ux���p0��E��c�gNsy�/x��W�!,Ixʬ�s{Ѽ<����`���t��w,ȬS�.t	c��pL`����e���_�+�����Y��ML��G��Y�����-/��N]��q�m,��JO
�\�%q҉e����I����Ю�2�J����i�UͱJ %s<�f�3-���8�"q.קuON�������M�e��_d�&��uqVݷ�X�Q�sw�����۹��A����`Z�'���wB��e�����T[��e"�_�֜���zJ+�������]ǒ3�N���%��=��L��F�R,��ѯb�6`�^��[�ɗ����D������Gv'u4�B��֒������X�9CWk�hǔtg�rso���E���~5������)Sl��������xʭ�����6'*�W��}��B>�8I�/X���S������K����Z�~����ɂ����S�N�ؤ<hE���"6���c8�G>a8ٙ�uuCe�x��na+�uy�����(��S�ǎk��<�&$�hM��L���q�:h����i:�� E��_�jkKܸ*���µ�%��#�|{5y/�?2&�ٙ?a녏У�S.^츌^�_��\D�^�2���=����g�)8c�Ӗ��t:^[��u�r�Y��@��E^L��u���}��>�gV3�S�����_.u����P�2�a�
h���$�Ν�Z��\ܭ����~
����_#�����B��$�bh�D��>���t���dÆ! Ъ��=WA�E�ax��Y�r�>v0�kq�k�ۺ����1OX��e�.�t+^T���TVJԬBa<X�vx���:+��1UK� �j���?w� ��"��7&3^Z����@S���>t3��i4�m��)UfZ|�WMu�GMR$5HEx���d:3��, ��ѡd�D5��gN���BP[�:��A�us��g��j��~�B�ʘ�I0��)B���nE�_1	9�|�vl��J�~ib�o�$����;0Az� �ށ�):�p@ӟz�%�S�i������A�q)-a��Vf��Kc�a{ᰞ�8P�^��[����R�z�"#��='G��Pq��J)�j
A'�	fP)��e��͛�7]9X2F�}���t��a(��b
&8��u4*B����ݟP�"V4�r�Q��?OF�� ƛ]���S�s��`��&�F�
��Dw��x���g��i����@Am�Z� ����QF�!�{�{��a���~��`�"S���0�z��B}��z���l�*.�ǟj�����R����FvT�^��A���V��bD^�..�Ŗv{!�[|��uW�3�����Y���Ǧ����k�a{��IC�^�הջ�}Z�,7��	i<�_���b�%Y��"OݝU���E�_ޏk�>5��ۯ�;\�����g'<hV|d1B��;9��=#Ŏ�^Rd��WsQ�{�p׃YU@��pQ�1�2*oO�D��)?�;�7˚+lE�����
�ly�(�8��h�&j�C.�!�6�@��Ɖ�gq�repB�}���Wb��'�����g��
gf+�3)~��9��]��{S.]'i��-��?p�5���ҹ��8�|�L�
iӻ��m��Q��_��ֱ/u��bu���e3�3�g�6?WS���r��62�$e|8k!~�pꧼ�Oe����JE���Q�F7����::�c���V�嵕�֠��E�o^�ʸr�.[����a$*�gC���SL��x�`?�PmBA?��5"�U�N,�E_�]"~E/��%^-h�/�O>:3Ka
x<ƌ�I��.h6=se��*�X
ͭ�9�,;�?����
��Ǩ�2gaҿvS|�x�멍8={.Hٽ�ܖa�y�Dwp��wY�F�e:&r�R����V����H|uS�J��ts�Cpy�ߏ�'1測2��H��z���a[?��[{3�[+wn�]��%��/Z�;s�Φ{p,5�)n�!x�S�k�����v}1�+0��#e���I�UA�=���f�����:��g�<5;;[�!��s#��£�=�I�\j��X����9`zLVc��D�8QvŦ����X���n�k�:;ޏO�&SDq�����a�G�>
����K�:�XoL-9W�9-�,Ӻ'�3�t|pԭ4��������v�/+�->ϒr	����� fq�^�������<趆7�M�0,�Bj��=o$8��W�O~,T��E��a���w���UE�po>�h�&Ĝ���7b�Qt�n��c�^�ԅ ���Y�k|s�I޷����wQ�����⹖KR��ϐ|�$(F��l�.�<Y�=C-�߳TL֧�3�`�.U+r4:%G�l4�Ot'�H}��|�
]��n`�������[Q!W��Mxg��U�W2���������q$_<`��0ߚ�ӂlä��+�N�Fny�<�V=z<��!�M��e$����_Iꬉś�t�%��Dqt���+��HH�gT�q�ގ 髡&l��?��&.1�Ju�'�^���s˭�_�
�&��N�cj�eP;�+��o�M�m&1t>gR���,[>�N���q��c���{�G1/�
v	x�������������1/��l(�3�1#"�9�D�����#���ʑĉѨ��ԕۗ	�9��V�΀�jf8�)���C�Eeg�)�.���)���Е=G��2�4aA.��<�������T% ��%���sS:�p�~@R��4�m��N�"NB^���HD����k����$"]*�FzX��3�T�k\|�]�D��6_����hk9�[o�wf��\pś̲1��&Q��`�=��#eo\�NA��:�|��U��rq��F����0���#���T+����p�0�0pʕ-��
��!a+E�=~Č
1�*ĹEH�Z�6�bP\C �1B������