XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���v��]��+_�Uލc`�~To75�a'�>0�m⿏u���M�k!C�.�%|Ծ�V��d‴ŧ�C52iXq�CQ��SS����m�|���ާ��U�v�-q���+����7(���YԪ3Zf�L��?ec����P8 ��]�Sr���xC�y��\8=�LRפR0&(�`��D���������g�S\V�_��������&^�݋N4�瘶$Ȇ`��X3ƴzEV
��h*B!���f8����K%G��_���&n�2�������H��Lu����5�@�c-�.5yj��O"H�9��E���̃z�u��4��O�
6W�����[:y����Ө��l�,�B���I�=�1�X��spHT��3��a��O�W���;����}�gW�A>\�i!mf������_P��D:��D���6��ILB���pQ���x��ƠӚ���?\�Z��_��Aw��f�k����P>��Y�)�0��%&[��߿?4_}��U-UD��cdL~5WGDY˃
�sDE3���i�x�]��;��#scUH&��h���*ԱUׂK���R�
����m����J�I�2w�[�dr�c^)�2Ѷ�<�����7ǳji.�j(<�豺.%S�JO�)>�ak~�� ��G�Z[��[��` �.v{��p V+M��@N6�ܓ�w2�/Ҽ�w,�)�N6XFL>�iE�p�6���N3���3��H���@{ �m2pI���c���aodV�8���~RXlxVHYEB    162c     850W��Ȗ��5��:�>��Ţ��xjS�,1��K%��]A�h$����uyt���Y�6?<}���|�1�e��"�b����K]/_����"���p���
���q㌅��Efe	�����u+��gއ4�t���g�~
k]�dҒ�&N��-��&�o�$����V���pӦ�?�M�Ӕ	��^��i_@[]��F`������
S�'�z�?ћ��a����ˤ�T�fϫ�iO1�N����K+�\���|��9Ĥ�0����H�h(>Kƙo�N
����t����t����1J`nX�`�b«��@4���e��A���!��<Cj�f��/��7�u	Oq&����)�x�'�2z��V	��A��I�����F�x�ZX��C����=�j�U��F荊[�C��7�A�`61�]9T.ö�y4X����.�Ku}A�Co�ߴ�)�`Ja�����q�=Z�eL����Ȍ�~���ɒ�d�����-6��r�~�̌L(�[�o�%�ޑLM�o�^��L��>bEbs<��$C�~AH�l?.`�"��GP�?�#hq�2F�ߨ�z`�a��� ��F7|��o��ҹ��:������2E[��2YF����3>P����C!E�w�����:'�\��j>q)�����_)9q\^������vǹ�x�#=�i��}�*�U��t�؅�, :Ճ��N	8�+�Z]I3�����~pC��D�*+C��׎m�Ut�s�Μ�|�K{�O5_�~ű!#����y�d��������e��/Т�͢��_�L`�c�̓��4:�%T	�{jӝԉ��8���c�:�ST�k�Û1$LDڞ�<I76m����X�![�׽��֞B��1�|7�x����$��f*�|����?��s�.d�.�|�P0S����
�f L�)
�^Q2�ze���=�ac���<7��|7B`�p�f�p����Gr��p���J�s�AqTl%	�:��O�������)I��:Y���V�/�i�{6��έ䊋�F��7$ÝF]6;ʮl&4*��h>I����nOzqmV!�4�(m�;5�\��#F�\W9���H60�8��?wY���mef6���gk8Jo���_��&��;���&I�,�"\��i����\��f���8�ҟ��{���5�������$CJ�<����F���w�A�Q���s�}V����$\M]���c:7�.�N�.󔦯��DE�fp$@�r*$�8kf21��ũ@<1�{g\�Kh�����Fu�G?�􋪧���&�RM���@�� ����uD#��+R�+Σ1�9m)L�G(���|:�?����ퟢE-�i������Ĉ�����&x���<�����Olz�7wnK�����ni�����J��|`e�+����й���{DP<�S�����ջѴ�g��d�`�0Ï�D���:�W�0��-���D��&�i��i+��by�bMK�FB׀�AU�Z���C9k�@z��,
'�	|���:
q�{�G8l�/��~�i�]�zQ����qcp�kCJ�r�����{\�C�z�V<F������vn�Ef���L��&��+���ڱ���S!��1��0#]�����w}("d�C��q�_����9�/o�iE�v*���i��e�*�̈́3�Z^��L���Z��,A��[@��Ys��`�*3hRe����9�Ju�/Ǐ ��
(Q�V�Q�ڛ�����I/wݨɳ���c�O|mК�I�OV������͋7 c<�%V*S�cMwtgR��(ȯ�,�����\P�χ�� ���y���#�0c@X��C��Z�K#��V:��� ��\���:^���x��z
�gR��͌)����n.r&)j'���pd���D�	 �vD�F�#�s����\�P�NWGW7��@\����|��� K;�Z�v�Y��}g�˺fk�25��B������32s�~..p���F6�ۓEe�v�[��HD\V�[�P}�>��=k��Y��+}���q^��;�Հ��S �l�,;�����q<��_���O�x0���,�+��7�9�����|��g�&