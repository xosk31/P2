XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����%�׮p�Ο
1I�=2r{&~sǅ����C�R�`4^��3x� �����y_��o�=HJ��yZ��#5�&D(�xc����?O"�'��z[~�s�> ��'�ŏ52U�u7�g��lY	?��x| �a]�t�^��(G��!Um��,{��+2�� ��K�S���){���	|ʍ������$����,^a�Q��:GCe�����N�XS����5��^��MH���8����4�wBc���;�ͅ^9ή�����T�s��=��4RsmԻOJ�	�)��>�X�0����!��#�5�V��6�o|�]C������&Zui���fT�Y��T��W�DE .4�u�uU;����d3+(�$l����b[�+WOW����J����9��=�����k�A>�B%e��Okl� q�J���B騑@��,�y�ݣ�4��� Y,W��W>K}���&;U�26F�t:�sN���!�p2o�e0�*�%W�fǷj�&B������X3�[R��-�1]��o���>���i_���>��5W�d�|(��O����n�ڦG�`:�; �M�y`���[��ɲ��[�� � �lP��eO�!6�E� ��� ��ObyC./I����UQ6����w c���6��&]Ɵ��)O��,���oJU҈��&!�9�S�dfcS�C�����Vr�"c�^2KF>��	T�<��ۥƹu9j���T8����\*n�A��
 *��,Q#����>{XlxVHYEB    5df6    1510sLn��E�37���g��,�s���G�G1���� M^EǤ�۵�GUo��ۏ�����lzW�k�� �C��5V��;�v}JgY��!Q�+���V��:#HQ�5oeM���r�.���E���J[�b^�O?����k�f�M4K������H�4���8d�,k�STH�͕�}ig+]����#P�u �"r�捁�n��Ǵ�gKb_����adm�Z4���2�F�Zp�nT��[�O(��&Ϝܪ�-����j�Ё��3�f��N���V�I�r�y"��$X� �郬@b 3���H�E8�	�[�!RzD�J����R$��7<*-���VX��l�(�����߰:+X��I�`1 � ����!�$��:�C1�l���֔�ú2���9+f��?��x�mfQ0���^SuX�0��]+��h�ߘ��`i���%OC�x�il륬�'_��H(��k��؎��M��f�,���qq��m ڣY��7�8'���s�`>aY����}ĺ�s�'�b��N(A�;װ�s�9�OO���u���RE�5xgPp�%l�5��Z��8�O`^����Gy����C?������ś�J����,̆����mͿ� y!��ɷ��@Wr}�����2�#�+�ld9Q����H�����<�I��(I!�P��T�i�o7g�	����h�}��J�9�v>[��:W�h�c4R�"MP��ԑ�p0�bĥ~��GS�)����)0��*}�^��_;-���W�U�n��VV�洬��JQ��Yk�0>au-�Q�W�	��Q��t|U���2fkt�-9���s�m�D����q�o�A����vn{QǮ��h�Um3��������?����D�ūA7#�����9�ڳ){�ƵG��Sv��f
UD�y��J�+W��ū!���F0�Kx��}/�����e�����0]�ńaW���g����DW����}5�'#�a�&v�����"A �/�����~���?��'FR�����W��/f�.�&��Kǝ丰E�UZ%䅴b2�R�m�_:'��]��?rm�#qS���궏?�Q����L��pj�:�x7�b�{�|+q�'+� ���W�*�ɓz�q�2}��j85c�F�v��}i[{2��/�p�Ou�t��������m�kU�̵�6fM`���X8
��Q�z[ے�\�k�� ��L�^���V���5x�e˵;jf�������y,<�u�Y�O(���o^ �%1�Ƨ۷[���,X��hc���3����]�2�J�ٟ	��5>���d+��T*�)"���)��!53�{;ޖ��|���\'[	��\��� �UkJ�"h�����X�����	P%6G��:�r���p��g
��[d�7�K��� ؙV���::3�F�P򳄫�5���?�����Ċ���=y�!}"�o���|+2���{�#Ӿ䛜S����i{���!�|�"j�G��\l1�E@Е����]@��n��(B#�1�H��)0<&��L%���L�?�X�i�0_��_�a���-�Qd:T�`�/ �ͤ	iŸ�d2�ia�׸L��y(���uf(�wQ�rYZ4�}���a�EӘK""�����(5��ӷ�^4������~O���ofz��G˵��ƀ���6:<��1����C��V���}��u��f�o��`�L���9J}��8�."i���vɆ�k����:�e9;�~4ӆ��$a���l+2���5qp�$�>��	K���I0��p�!J��I��� ���k*��˞� ��~uٯ���f��C�P�*���_V(��:�ǥ��;�T��F�*�_���_�>��l�~oL��ʖ��0���sH8�p�%�z²&�\p�Uk�(�%[���wqT������f�@��n�v�&"�{R,�3	��I֛�C���	�G�\������О��S2=ѣ�'=�Wӗ���ɪ�m��\^���Wr�Br��)�{\����y�s4Ы���/������
Bur٣R:� ;H�_X�P0� �_8�=�ћLo\�y�h�Q��
��Út���D�^�#�M�X���^���n
��	�����Oѓ."6H"/Fq��5�?���6W���X�ɇF(�mJ+����\��v��B��F���ο����;Ѷ���Mbw(�޹�)V�'�^*��tn���{^��|���G���ȥ,n&�I>x���z�
�?��TW��dyn��F���͋�{� ��8���mP��PO�'����R�G&
J�(%�j#{�W�?�v�,����R�v$?p�)ٞ�b��{�fl�;KJ=�%���nH�ox��F��%��
��'�V5�+~t߷�o$� ��pm��LSk�(���5r����Y�[\g$dg%���\[�u-�F�\� Lb�����ʏ���Okө��g�y	i008=�J�C�`�o��]�Ȟ86���˂[��a1��櫧2zVu˛��}kf	N�PO6�˖����q_��Z��_z߾x���������=���~M���l�7[�q	7���Ed� �=C��vc��B6�Y��I�l�2���F������J�|@�M=�F�/W�K�R����Y�q1��&����,���(��	�l�_�1�����j6�E���y¨LT��g�?�z5��� D7��P�S'����2�.%H�(��W��%���q�����JiI�XDj�+-�Hh�������3�J���@�	�ٳ���`]�?�aiϜ��3xN�ة�R8;�*�G����ky������ji"!��z:��uf,�>��獻�G�'w7i�����r�@YB�,1i�����W2+d�e�&t{�Rr��=�1ác-���_�k�A�E]߲��R7(��Kcrw�� ��ؗ�g�7������1e�K��_e�"��ob � �ekkԚ�Y�9�İp��CU���l[}���^�W	�D�P#(�u_f�eX������t]���qt�}��NO��1>��*h>=[N�y"��%�ت�u:�)����A��:�*r�;q0�k�J3�YKi�#̶.�/۶���e��f>���?��$F�
#���I���8<�$�Cؠ 6��\�*'�U��ix*���KgAZd=���w��ܲI��t�g�¶��¹���4N�y��kO�ȟv�-���z�̣F�-۰�9�^�yu��J7�?�O�ݼ�Ԍ�oՆz�ԋ�`^�}�"�����bQ�W�f�wfFx>3�o�7�ͫ��1�G��
9�ɘM���y^��MV���=J-5�c>i�O��i۷L2�b���6�&�iYэ9�ӓg_K�E%$< F� �3�Y�H�����Ņ��ӊ�Jϩ_5{�6�_�9*��1�Ҵ���CMI���p�:駉�i�Sx���8��2(@�o��\w8��5?3�2�����{�@o�v����v��n�GW��z[��Sy�C[�8f��4q�����`҆��L�4�l[�}�t�X�5ŷÜ�[
�-"�"�O>Gi@���x�B�C��H��H>��û�9Yj���4
9=Vi��^���^pƧ?�V�z�V#\^���,9m�����u��̥���ޜ�㘞�{�,�#��.�d�{�B+0mv���,�C�I�1i4���H�(�S\IZkي��ʷ��<y����(���θON�n�D�)4�9�'��[�G ^ٵ��0$��t�p����գV�����\̇ch�F":FS߻�yD���r���y�z�8T޹��Wc��.	��5E�JA�X��GUlB���z�	]��<�)<4xr�G���,�mo��Մp��u'4�gʋm{�e��w����d׸ �@Fz�͑��-<V�0�\�c9D�y妏8?Ğ�`��/��(��wl�n<|��\����a6 ��YnRHf��#�Eyk��#���hz��6}�w'mi��ݹ�.K,�ޚ�F��ӡ��m�"bH�|�~�����
Nf��ʏ�k�o�Gaj�����+�8E$ұ� �k�F"K�{�fC�l�)K婞�|Th�������b�!��Y�`���Y�m���������8h�V N)۫褯~ɓH�ͪh�}o�g�J��;�������tƭ{|$��z� k�a?��#��kv{�Wig�0tR���h�x�r:�T�|U�F04�8�
��љh�}�W�Y�+m�1:��gԱ�y7X����Hc��`����cXI�K#�����l�g�(�F�I�荗�VF��f=$_���ɲ|�dk�j�c��0��>6�H���t)i�F�$2�o��}���5�4�4䕸&�dS ����H�[��{�DȵT-��W�{=�хH���� C���B���(�Coԉy�WQ9���^MmŘ�2���+3&�r>��N�Ȁ=؃;�uΓW�OW��2:z|\��GMl�g��:K��WmDd��1A��&��L�u
�S��6A����KU^-���4E�6��ow9�M�P��Z!��A�0\8�ty.s��]��e��ඦLlC��{4�KT��AjO�:������ߋ�����Wr���20yy�Y�~&�S�(�f���Á	��x��Ú)~�g�q'V"^�"��Z^��Y���"�S0�1�N��#1v�C�C>6쵘z{���Z�bN�[��㲰(,9����A�&��ꍿM�b�����N*���8�%j�㝳�����5)��q��7�u~9Lc8NZQ���rv �s�#E�\/2~P��XTϕM
��绻�$Mˤ�U�y�Y����Z�\��y�[�P�R��y�FGb��&e����d�$&�ǂ�#B���n���`1����M�c�֙L�eg��K�����L*��"�@�h7��9�����]~v��	���?�b%i5�,��LV����{���X[�/7�$>�3
) R"�1
z�����y5�-�%&��}r�������8���%63=���o::ڡT%����{�6;�O�<M]�0��T�k (O�FT�@~?�[1Ee�2�c��x�GZd�z��~��5�Iy^k��9�\1���Fys���Gl��|��u���_��Nd��M38T�q�Q͘dC�h���N8_�V׉�p!|�>�0�)�T'�S=r�I����W�!��G�`�ȡ.~F���fɜ 9��Ў���3|���(Yr�ߕĂ�߯� %@�Y?��=ܛA'�/�/y�
瓦N�t�O���BAc�����"ި8;���u_��	;�
����  ϡ�u)�`dT��4