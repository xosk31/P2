XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��p��w��"�Pc o_���U֙b�(���gк[F�;}8'�x�9�|�$ըU�&��K��S�\>췢�f�������n��ĽrW@����3JT��cY�!8��ez��ȧ��1yL���!�
c�&0�*CL\���-�%�za�������1�Ř84��2�Q$�9�����~��a�jB�[FD�� �ǒ�!�)�i~!GA����=P^$�=gY�|� ��!>'�:�<�� R�0%UB�0�Fv�ʏ��q %�o�t��S�D�6�����x�礤���\�٤0�3,iuE�D�"J�{�=�iC�<�ؚ��/�TM�zу��mQㅬ�C<�i��I\);SL�JW�
v�гh�~ T��7���-�K��[�k��t@���Ig��
�b�]��*5A�@�W�U��1�%M"j.5�@*�X�\X��SK������4W������ۿ��RPe�c� �R��u$�hGؖJ�K,��*�q"�`Il��
�������g|:x �X�b���B��։�Ƌ��M ����+�i���_?3GA3^HBA� 	��%�p�ʿ8����ƃ���2�_�ʱ�k�=-��x?f<D�9S��<2�1f^�Jx�x�/e��@5
�C����s�����-��L�d�\�Y�)�I���?��5��;�;l�0�V�c�t��_&�\��h/�P��8�\䀏��q4���/�8�oo��a��\��0{��I||$M�XlxVHYEB    32e2     b70���`�*�[���y@���ZjGar�3j���Y:��q�㎑�2��ŶZ�(��`��n;�=[$�t�z�5'���燔�U��Ɍ>帹���b�>y���ȠC���a/��/9�`w�Ҡ�ZB]��>w
�$� ���{o�]�?�����s�Z�&W�I���ô����m/y�����)ɢ��d�<�ΞN�6	�41�yv��C}��i�M�/�no�L�O1{�:25/'��]ZE���ɨ��]��_D�'C�>������qtDY�m��0�Y��k��C�B&�D�z�p��;6��nYP��)�_��jc�RVG�^,C�)��m�B�}�Sթq�GY��&?�Z~ 8��Ԃ
mV��;�{�nr���"�6~�������z5���;��/���2\_`��ꚟ֠��7YMJժSn}V��&�B�+�ۆ���u4�,�BkG3^��Ĭ���X={*��E�k�����o#
Z��rJJ�p����Vb i��FG���2��,#��	D";�D}�G�������~C�&����_*����5�fbs�$�/8販w�a�a�W!Q�#�`�g�o�z��	��5N��J�Ӽ������1�<�(�����I�Gג�!+�<�R�MR���y�wD�,A@��f=\X���ѳ���ZN�}�W\�@|��UW-�"1�U��ɵ�~�a]��ϴw�'�~"�'���O�@��{oߘ~ܥM`0"c����W4�LP(e� ?�53N��V����4^������Q�mD�o<�|�2G���m_��i�H3��%$�|QŪ�=E��bA��O1N������]����Ҕ���:�g�����r?��	OWY�X&������$�4/I�2��Y������@�R����|�J�V:|SS#��ֽ�HJ.�� J|����ϝ��ޓ�b�{8Gà��A��ʎy�ز���O�YNQT�c�)���e�kEͬ�DD�n6����k�:�����R*�s-@�	��Yltr
Ƕ�Ҁ�W>a�����0�v�'���S�ZM��|�Z�0]?���؇W՜������a
A�=�D�S���`ߏ����ֺ��faj�2�ؑ���\	���4��) �2���>F��`��4V�A�G-��#FVמ�e�F��"�-��M}(�;W��<.Uk�j����BB�"����$SbFR����7��?�#��u7e��M�z`7��#��|���?��lD�xw�/ߺ�佮È�L��A��������L���rh=^�4h�p���u�"�?=U��Ғ�M�c&n�V��Så�g?F��X��A�U�6�h�m��:vB��T�kA=�ʰ��4K8zy�_Uma^��.�]Cyo�	8�eB����P�R���ʸ���2P1q!�1��Bѧ���讹kD�}���z���D�YP�x�rH�y�G�l�f��+�Se-�fZ�mąZUx{�\zp+��
������8s�����7�Pi�]�;JD�^�t�x�:)��!�@�����g����{�$�/D�\fJgDƃ�@_��l9��t��Ko�E����1����	 �Wtmr.��2��ՋU!�s����	��γVF��%��N m�rW���)6���_.L��H�M=v�V����aA��ڎ�H������O��%6�l�NݖNQ~�a��g��h7��W�n��p]���
���
�6a�ym�em[9-ವ-�e
�ev��,��2rd�����`[�y���vv㒪78�����]W8��n������C��z,������F7}�)��<������k�F�M�����=\~���i��󷇗q���G�X/
��L]|�39jm|�G���qM�D+�F!�6x��B[-)�22�����*q%F�D\�׎� �ޖn�9�ʧ1
~�bV$;�nhS��.�!�6������&e㿷M�J����4nW~�6H�)���\�9o'E�j�+ڰ������ݰ��K�����B�� @{�p��4��oǖ+1�k�������y��SƉs8KbD����Dt[��V����qQ�	�=;x��T�&'��4�֬�wW��=��Xp7(�]Y�H�/��N�9c��I~�P�����7'lª{�Q�M����/��^a���A�B7f�҆�3�sU��^C((^�Zi?~��ѯ������ ,��Go5�2zj�J5�o�ӊ�8O�
z!��^����CC�DZT���V&	a^�?�Uܸ��wH�_��X̱^�mג�)�S�-�=k� d-O�v�*,�������6+Zi�G��C�Vk�!(ƾkڟ��JIY�jS��'�5ge��#nϹrV�x������|8k��q�l:?���d�5+	��*ř���0��m�AM�X�Ԙ9}�v���]+8cA�VȃQ������{�Ԁ.;�Y5��+�b���ޢ�9U|i���Ёm%�5���g�-2c���g&J��Oe��s����и�Ƀ~j`X,W���\��!�J�Jʥ"��_ ����7��b����	��i��C�	�k��f�f��B߁�ɕL_��`�.Q�w�Jh:a3�K֔|�R��T\~�j�CNt9{x�@��H��\8Ӯ��$��|��,N&�e��M�$�r����.,���4�-m��Zg���%��XN\{y��:��Yq��!�95�J��P�x�Bͩ�0��2�tMo��#)�5������R.�q�����������Spm�Νݼ�@��c0x upH>�j*~�t�R1��|��=�eU���}���������"���)�6��:�g�I��B��Y6�svשEiCRh��;�rF��o�{�A���U