XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���*�j���~K	^O�R�X݂��C^���+L������:� D��'�_��F�DeG	���J����%�x+��h���?�C��ŞB���V���H?�f���#�����B�N��2qR���l���{8*!�X���F���`Q^ײ�����?P���_��N��>�z���V��"�$��!{f�������A����P��ܝSjzK%�6aZ�O�-�
�z.(�Â��g"(�aȉ�+�1�tšbD��O����E���I4ͮW�bTYZ�,+�y3{!p��.�4o�� ��PGEG�YVdyVv�-g�<.՛�K+/�sd�1�m ������14����C�#*�XF(M�:�M�Xvu����?�7�yS��5N
j0�5MB�n'�-ի��1(�p�/�E���? �.�&��<�[�.C��<��^oµK�E1;?|(@=��Í��͡��	���N��!�������\q�U���E�2|ҝ�u��Dk�6���в����c�)�O�����m��M3�^�b��<�zX�P�=)3��m]Ţ(�D��}��«|��0V�7��8I�ơ��w�#�9�9�n�dv9�&�E�w�Ҁ�%��ݍHH�^/F��̅�|��������ς�b+��Yugv�_�(�� �X�݃l�7���-DIQ,���x�C����QQV�K��;DK�o��J�)ę�,�vC᏷�J{��9��웣�XlxVHYEB    c6d9    25d0�ǹ�(��<�����ߔ]N^%
�l��Bp?ƟrL�����I��:&�	F�GB��n��60\i��g�{Ҧ����b��.�
5�t�&��#$�3y��OJl��
��0JZf����:��e�(0�;q�	ҵ�Z�c�W��:d���.���z�9�Nץ�J�Ip*���Ȝ+��o��{��d"[A6oVP���Ab>�u��u����5 m�R��'7gX=t�x�sH�3���J������֑���)����]E�y �Fj�yԩD������h�O*��e��K"�K�#	�.���Y#G�y֞��#��Ÿ�	��{�-�	������L݂������d���c�L����v�⒮�����;fqQcZ���0���J-���Й�1�5Ƕ���^{@;<vrgm!7-V�f�מ^��{�T,�\J��C㙌�&��\v�?o����-G6C^h6͞�V=&�a�Ha�:�a�Q~�E����>a\e>|ܼ<e5�������|��Gh!����C�n�����Hp��;�f+%�v����#8O<؊���l�YA].�߇ԫ�"���07Gz%YM)��wy��sµ>zt�eb	,����Nؠ}�+�O�|�	���[��.��>ل,O���U�yvU���{as��`	���q�:��AX�͜#D� ���s�-@��/�Ӄa��A� e�zF��Ə۬'�,����	�-O�yr,[j^���?~�E��_t��r�\��l�	>eP��6�U��x�����n���i���ڶ�#�\c��^D_z��%�����\�C8�mw����E.* A���<��f=�CEcX��W�l��l�l�����@v@�3�ڔ�̐��n���5�f󌣳jށpM�c0�^�9�t�Td8A��uI.�D,���iq��7s��P��n�>A����������9�m�V�[��bי�]0d�cw���Ċ���0d��Se< 	�;2	���k��d(C�%�沟�բ���-�i�ل˾퇀���q[����;?z{i�j��Լ����9ԋ���^&YN��4S��y[lb���tm2ܷ��f�s���/��_{n��(�01��I�0��.��w�H.�e =���B���C�A�phV{��=s� 岗K#���E�ށ0 T�k7��g�(�4BC���Cu��l��1�>@d�W�p�J�	�|��)��r���v�;��4���*ɍ̣{���o��a���o�o"���[��n� ړ�_�Jaw��9��Y��%��6�CO�㄁e2����$L7l�cW�$Yi��:��V?�eSH�qݛ�o��_�V��"/���ncӫ��o�wyG��I�q<lб��5��b�$Fz��<����p-�4��ش��Y���e�Od�Y�b�Yv��j��
a]���S��e7jO��!{��<�5��:h��_QOd־�em���x��1�W���	�N5��ko�;�O��pf����6.�)�d�:��é�6��'��=��ո�@��'�}��sZ0�BO5���O�<�,���_�rv{�+��_�0"lq-��jK4�n(Cĭ����J���Z�ɉ��]L���r�K�'���PLt=[�_�0I�o��f�bt�T�M���&t�*�CP�L�ѕW�� t�|Y4 �;������p�[����)?�i����u�1D4�	���޺�=�|�
��<ZR�`��I�'�������S���)���v�I"�{MHx������c����E"�5ƴA*��
L��S)�i��gF�a�-�y:_��F�%s`Z�����y��M0o�l�q'��}]̈����?��$�6���n{YF �l\$a�� ���	n5W�|��\&���+�ce�~��������9���7�����:=E�[ۗ�Y�v�[�}Z){6̞�k��;؋k��||E)���\6��jm�N_��틼�#�fng�� 3R�b`����&ƖD����l�mɚ2�y�QD�v��B�� {�C�Zir"lQ���\��8�K��(�-@�Y�a����E��>\��+�J�RI���=�|�+ŏ�����z�c��^�w��9��`����+�\���֡���� ��wػ��J���G'�C�z��ȷ�T�(k��R;�PC�f�G���S�╡z+�Z�F9���E˸w辝M�m^`f�_�w�{K����T�n�C�L�:��^Z_b."�7Զ�ڴ�Ea�̟������Ȉ��6�{������Ɔ��b�����!p��1U�d�z+�N���D��d�P�z@3�{�a4�n���Vq�;  ��V�>�\���[��d�����X�f��_5_�%.�q�|p�'�7�^�;��-���e3(���ۤ�(L��ƚ*����+(��wL�ɛ/�M0C�T�z9���V�y���)7?�Y��ۄ1V�]2z�<�M�j�4�!�I���gP���H[n����S�&9�Y�,-����� ֶ�,1n�2W�tDK�S^|�8�:�p\�UmYI�u���C$��Dc�P�,�:2 (�ǭ�5C�v���ѽ�m���=+��=ba�(o$��\���'����`�~�istY�]�MtsR@#��
L���ZG�f�TWέ�w?(R|��x�=CF6�j�D#���g��c��>OI̦#��or�_��|:$�jnN��e㑳C�K~��W�J������8����E>��SKH�sL���;��fZֹ,���!�Uo�o�k!͞���ˢ�
�O�w�R��S��Ɇ˱����[J�1�OYWӶ������l_�v�>���*�Ω�0w���{r$ы�e����,�C���7����*,ip񯝖�yR���(	��Ig,~�ު˅d�����0�l���(@��{%������Pu�9H��>��.�V�M�5�d�_{�>��	+9E�(�83�p'S��6Ƕ���5UcTfF{ˆ�/�w���}�(��Y�p���:��˜�O�}1:�С�0�(t��EkXy�b�3�<�/��x�^1t��hŃ�y?z��3j5���;h���'	��F�ݧ2�"sM���g��*11y�O�z�[uv2A8V�N�&�ig�����n~Ajܥ
{�1|ˢ�ǻPr�I�����==����������#�l+7�&��<���|�z��D���8��茶�$Q���7�{���Kؽ��5�x�ny��QK��%=h��Xjv�]b5���,�JG�/���r��P�����L������^����[j��=�3���q�����ןb4�L�<{��|�6����[�!%I�?JS"Q��������Gg{��^v 0>6I�d6��N:f���t�:�N��U���â�0�J�mS��9���
פ�?=�BM�M�ݞ������c,�����zœ��Za�#��g�p�|/�)���O$A6��^�y&�
�8�����&�O��W����n��tZa5�tn�Jڧ�qA�\Wi�t��#�I�/���.O�ߪ�Z+���^�}8శ�-s�b���l�����(g��)/8�6��ȑ\y��N��唚��i'���IT",H��E�9|�]
ń�)!���ͷɞ�n!�⿿�{�"��W�����'-����Q2��;4)od1����ߕ͠���i ������}0HCn�X��(�¦�pt��K4�ܮ�S8"켪�������A�@�&b�X��MW[95��9��	��Y��*7�-��8F^�������ť3�+	%��`�H��ϡz���C�d���A>�,(4�J�m!g=��O��+~�Pm�u���e>������/�^������;���� 1FU&Ɍ�Q�[�ʾՑd��~��q�>Ԛ>��܁��$]�?ێw;��j:�bS']E�q�8�����$oDB�U��S���g�����op5��
��)VuG�ه^���z�SDj���r	.����N�a�>�~��>z9�c����#1�*���y|���o�X��8/O��>8-���,�R�zZuc�5'�T����{�kp��C��e\��*,y�{+�"$l3Ȟ�K��(#C��-�=��n �����|�Kv	>�S�Ԣ��0�B������0;�1���R�M��\����#���:��+����7�Fj�1�kv��� �I�W��o������(w�O��z���l��)�c1_�.�xR�����p�*l�����"+p�����ƴ��|��-r��6�p"B${�6���3j�1��2�oʕj��`���B�e��������Ч��OF��' [�G
��F@�Y���{�e�ǚ�N ��ux�<@�	�Ey��l��C\�(��D����e��F�U[b2DV�5���vJ�6��D�/�6����6_~ �S�&3��������d�q�A��g��Fr���=������cԷHbu��{�����xp�<�E-j?��Rw%�$}�-7VW	OY������]X���Q_�TQ��.�d�Ÿ|��%	�}�휣jW�'�b�L���?�m3�Ɖ�����7Zb]��p�C�|p4ұzC����n����$V/}�E��Q<�~$�%,"<2�Ė��x��¿��;�OS o�#X=��>�D�m�nܛ�O ��V�ş�K���>\��W��n�F��U5�ি��aq�6�3��\��sz��ҕ�Ќr�V�M��V*�(Ky��C�k�Po$`�T�X!_O0��f��Zl�,��s�St�ab�U7�"��~r�ic����5ԁ����v�8��ҩ�EW<���m�ʧn&E���P���(  !
�"�Kz��el�@��`��D�wW��h�t��\�X�+�XT�D�/��V���֛���SS�4UV���IS��!u/"��-7�s�ڐ�-��h�A6��LK��<M����:���^��)�#���t�QR�pPH�d}�.d�$	~ioB<����ZHlCܫ\�;g'�9f�3O�7I�\��Fh�,�8�q &�~['�����%ȃE��[@ %�b��;��+��0[�٤��=	۩�r�B<��Nz�YT��!�^Ku�} M�����4�o	��F�ɢ��TPJ��@��k��_nt�y+ɞbD�`п����ϑ�9�3�;:W��\S�?���6i�����Z�@�L�M��읹��{���b�C��w�� ���$<�%�͢�
̀��?o�/��ڷ��K@��\�� k�L�@�����L��J٩	��Bꐝ%��:ڸ�&OϠ�nC7ە�.�,qw)_0�.�}ZOT,��D��)P�G�  ���?R:-c�۹֠]�D��X���ڵ-��f9]@�f���{Rf_m�nT>��t� ���`����l|˶�`׿ĬH������܈��_��z?�Xv�5GTn��u�j��e�S� ���+ݿ�!P!Ƹ����:>Oľ��W�g�]���&ZO�� ��UJ۠ģ�w��~=k�k�q��-�AM?k��y-�8�5k$C�7p<D���)m��]�Q�?[ �"=���z�U{D����>�����Pu����S�4��%G2���V���=��g�k�S�+��
��\"��7�0�c+=�K�*û>źX�M���,S\ys#�o`Y�\�c|��"3pxǁE�_O�
�����x R@���I@�HK\r1�Ү 鍢�vw�I��xR���Յm�3�b��4G�1�v>3[n���u��5�AI�~��|'���0i�_7:����jH%�/V�t������UH��.��I�xk�T��<'��ڳ��Y���~y�&ٳ��W:��� ��g�O!*9&2(��+	�F��9F%��zRh�������P/<녠�� ����"4i��O�c�n��is���0�*����<zJ�p�x������'�����W�d���5�Ƞ�e��n>����{R�9RNﳴ�t3����'�]#��n��\L�(��>ہ�	~�i���2\^?�ut��0CODsz�$H�Ö�KX����)�``���&�^�5��b���W;�!�r�P7�}�bQ��Y�Tv�(��6܄	.D(��y�\j�h�s9�r�܎�}o>�N�N�"��ݲ�򍉝�	������� |�[f�I�η�'��F��h1Qg ����<c�ّ��b
���%��<��%/�0g�>��������Uܚ�Ǖ�PhM��{�+�7[��N�9�qV�����@����%#L�]���^x��ډg��x��f��0j��bf�)$ppd�Ń܅�Jn�q/Q*�_��r-5x6��n9���	�L
{���9�c-}���{[m�ΰ�f�'���T�j{n�t���9_]����x�w1���Iՠ����R�I\�m�@~r;
�!�"��XV��n���C1��i���|/��������fnR2�`@\����W�4o.�;��_��6�
�w�<򼇵J�_�ދQ�q�����"'ۅ����v��?z)���
o��g�˄�m�H\'��[3c��Z�r���wС��a}S�vk�tt��뢋	!n?I��	Q@9��&��u�vX�V}���JpA!W�V�������~�,��'�T%�*q�qu�/��@�
 ��v��"*l�F��G�e]jሖ�:�j<,?�yH~A�
�h&*�rqקf᩹#���?��4��w��~����>���o�3�s��L	�ք$�����<0���-Hzzڀo�g�����ƶ�$?Gm�qϦ�=5-�2c�ϧ vӟ�}
�9p���TD��c4�y�c2I^Q�J��ǩfm��oE��d��W��]�Kv�˖��z�k���,� �I�H}/�hOa�#�Ӆ7�^p���p�2(+�Ԍ c4���5���_ޝԊ"V��x�%��Hd=�L (9��0C�jrs���m��
����7��O�� Lw�%����*)��U<��@.�ԍC��	���T��FU+�̫)w�@��R�VQ�(R�;��t�<W�ۚ�`�v��ֈZj�$g*W����=�rc>:���q��ANp��Y�vӈ$ռY��|������37�n��������"ʣ3���<G�F�Hxx�]T��-Vb�i����n��/�B��m�=���I�s�b�峳��GI��gc�"��a�{�P����=y�Q���K���fh����"�|�q����b��E'�Ӡ��Z�`���֭��;_���St����U�X90L��Nf={��b��8Ϲ�S�,���H1�,}�o>XC�P�������X9��V�;Z�V�<��Hʠ�ٚ�jp�x��������GlX�D�{���)������5����>�\�jU`0�O�^��2�ޜ����qsA��"m�c3)���.����+� ��	k/ԥg�>���J�6���-M/��-Ꮨn�.��7q�Q�D$��䩘�S��U�\���w���/��E�Vn�QU�θ�j7��@���h�m̾�j��Z��������]��e�q���]o�x=覨�J���L1w< ��f��PbO����<%Y3	���ۃ)�r���@��wk��\y=��Iwڰ$Q��`�Ӛq�QUp�0�!������.���`��,��#����ps���Q��XU��
��3����V��H�Y����?G�7r9Il����R���ZᰀNgx�վ��Z,4:�f���5�����z������Pn�A��%Sŧ�;�&TI�@�3��Xh�Xs��D��mUN���'��������΂E6��ɐ�1��Z0_��"���gv�.�{W�i-��S��㊨���j��Yn���V''���_�Y����#��qO��Z�p�"�}�7?��L��(8�e�������̌��(��[�%BV<����V����!��p4�Y��]Eb��U�RP��Z��꺏�X��?��kW�-M)����~���R32���� ���ӳ�P�:�ћa:صx�c�)l�Gr/�0��"�=C?"���U>��̶����[��(P��x �����C�hu@���@���?\�7�r�n��H�B��������$��qA�h�lh��s�;��"%����ʿ`�,��9�������vq����@FQ��&(��@�������Y����G��Ԝ�S�9�~J����o��-؇*��ѳ��y���^TE�ĭ7���P<��wH���Z�ԑS ��!����c����lW��7�����>ƶ	��,,Í/�2�hע����X��"ӁV����
r��djz�w���ԡ���x6�� wc�`�/vt�OA� �:nF�P��;Kb���I��8XM��'~�j���y=-4 ̮����?E��Ur��v��"d�#��WA���n����2�n�цL�������ݬD�%�7Կ�_��Qe�36�❽$ݣ�jQ+L��͢ś��L����VXQ^�r� \V�`�e��6YF,ߜ�EuX��膍�� x�sY��yf����9R�� ^=��U����'�x� �T��nO��wFb*RxTǶ�dv���2�+O��@�����29O�r�-#�<�V޹k��/�'憉T��bc2la��Ѹ�T�x�9������A���4��^����1�?b�t��Hp�Zu��q9��	ଂ3���
0�]�d!&�D�ui��9����Wl}��dzl��?�4�f�Q)OO�C�_�h,6<��rxV0U��Z߮+ق�l��Ѥ=NkGw�q�W]��Mf�LXļ%�csd��
8N	�οm����R�"�jP3^j����Ll���=�d`v�{I�ᦎ���5�;�{h�v���"ĺ��+[u�o�>�5�%�Gn��afMjD�����#b']��ڹ�<	���(�6[�5d��}vo�"M�7FO���k����T�c`��ZA�Y8/�_P��q��GEo $��!�uU�N��!�c���Ç���T@���1!�%ޤ���v�<��R�ǆ�zpG{_�+��4���@U.��4
7K��y��X@��3�nnVwFk�-���JSX)z���� +�k�L7��MG���
�$��TE���������p��!�)5'�'��3��Y5D�����d\Y`�M��M���%G�iԓ��ѫ��eE�XG2�N�N��r� |:�q� ��l'�ύ���E�f� ����P0��e��X�y�->�y�*<�I?)�ˠ��$�nw�1�}��l���H��\����'o�l�7:�جS���� y���@�i�V��K��R�X�B _�ട��Ja�"�k��x#��	��FU�T��%�`�K�iDJi��w����tb���&5�\trrN<��g�Ⱥ�
Mצ'C����8���]�&���^���5����Ԗx��n
5�i
Ӎ�*�Jɜ_������R���*H�23�K@A����H]�