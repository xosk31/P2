XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Nj\">�*�f�dNJ2��wܶ�B�cΗ�d�La�~ë�~V�ܣ��yt΅��a��y�b����l�� t�>�i�W��Q�,Qm^ylM��W|��G3�M��7��<W���G���Di�(T��6�F��V�S�>7C;_�Xb?�!�8�p�b�JZ�D��(H��,6�*����~!�6����q�r�Ϋ��K����z��Jy/@7Mt�8l�ü�6��LY6@N�Z�Aͻ�Ϭr�r�I��*���E<mDy�2��\
���ܗ�FJ��xu��E�%7�N���2��֡CE{��["/�>�ѫ���)E�I3� ���,�
��cΟ��:R��JAj�`=�0+7�z�ր���&8���$�0�����Y�u��Ӈ/��T�קąiW�yWDC�9�yQ��U�Ұ�@���DFn�H�'��Sf���-�愩B��d�-\��cU,�<]!��,wO��"�X?J�$�l���F��I�����s�H���!XYd"�(�Y������K�#�����v������i����D��!�x�7�}U��$��$�R�����=�}���@<ްǇ��籊�zXÈY��q�=��ـp�01�J������X���k��qB	�ˍ�#&�+��,���UE�Lc�ϥB�
�ͱ���}uMBF�;�j�`ߛA�o�o�k�E��[UTZf@D��;R��!��9��-�P��샸b}%�J̬|x��ɘ���l~4����0XlxVHYEB    5909    1550�qc�Ƞ	��k�烴z��-*��k�@FK���]��p �^=c�h{*�fIzȈ;��m� �W��i|����)y�h��N�%��o�Eh��j�Ψ&��XN�T� ���,}Ѫp�����f��L��3`O{l�樝3�tU;�%a�Sr(A�C�� ���9#�~a%��K��}�9�(��AUq���N	p��	������Ĉv�K�bh�kd�@f������OM�(��r~��H%?�?�G{�|1Y�SBBZ�B-�m�Lޭ�7�АC*|�
�hjjE�^�?H����"M����$[�L��؛���R66�֮�z�6oy�O�$f	FАհ�o�y�W���;>e��j�U)�{��]ÞN���{}A5���/_#-6�v	�5�+�GA`c�^�w�g���X}<GHd!��c�w�U�n�*�j��*N�"LB`�
^����V36�b��K`�q�|v�bE��f�Ν�e1OS-Z��XE�V+���%e08�(E׮X�E�*6�^?i����1��9�[�$��l�].iϹ��M����hh¥3�Zg).	��9tK9���p,�2�ꕜ\���0����P�v��J*��H �������ʝ����� �d
�)��bBf���r/�o{ۿX����<a`6��/�B�B�4,���7�.�L�ʵ�pfh��Ϟ�g뎨�j��1�-33�?>�[/��;c�x�8k�K�ԺX/S��\^�˶bݚ
����tI���Hj��of̓���\������I!�*�>Ǆ�}�w���C�F�:Q6���ʈ������G:O����'�8�wu��Ӵ��X�,���O��4�O�eC���m�C*�5���xF��S"� �9e�s?>��/��IW�Z:���67+�vވp�z����kjU�W�H=��J��F�6���K3J�7�e�>^��}��bnݶm��T� M���I�̜!�۲���Qř�J��܌`X���hG����lA�N�!8��]���$z���V�J����Ʋ�,��t|�
*��ka�Ҫ��6�FWejɓkS]ZJ
9�I���y�<R�C~�<������?�A{�2Z4����O�G�a�yS�Y�+U-������GJ�ky"ɧ##1ŷ���X��i��RG�+�G��n}-�k���q�t�!/%67�#��/�:�:�]� +h�#
d;TQ�l?����/-amXj03�hY�`H�2��� ݑԎE���܋��m���/&�z��/��4f�STE����c�bf��#
�����΍�F�1+/^��j[�E�
��t֬�l�S�+8�U��W�ؾ��rM=�H��s���=��~ȼ�XN��,��EJ�����O]p�G��3�A1*�F���AQ3�*��2R�w�i���?��;��7��	���D�1m�H*��6������}B�4�q��	�Cf����}1TΚ����3)�>v���hq������j�Z��d��Sj�p(��ԏuD�J���wطQ�ƚ*�b�7���X����B�@?&����5�6Vl��b�>
��,��̷@���f��<�yV0�����V���Uk��v��7���Z#/-�Ų�[�EҰt�1��������8�($���U��r�KI�2��?̅~�$���WȰ@��&�g���W3���J(���6�#��]_]�ڃ��7)�T+'<�������Qr�~3y���q�/�arʕ�ǵ������"���^���RUh�nK�o�F�����5��`�bV���H��o�#�|J�#�'(*G0�?j%WH�nb~�We�h�aB�:�����������"�-�vI�	�5��������H足�� ���R������}@��\��/<J��)P֋����`-s����hb(y�\a+��d�<)����5qk{�� ���8c�Kjȳ{V¥;г``Z�N�)(�X5I)���n���"���hsqP[���9X|A�{ޝ�Q_m4S#r>;ۇ`�"%q�F��[�e��[$�/R�F����1�"��ӰJ����_o͜_��Q�ܲ�wݳ���`�E�]�XLv��x��7��s��̴e�cNj�QAΧVg�AOU���Zx2��@�gL��=��@��&\�A6z~X� ��X���8�8F��xԢ��s_W�,€A8��a�@�h4��P;W49l<��CB$�Ց�jn�I��%�Ba�+Fel�Wy%m!m�^ E^c5ǫ�D:�:k@3�>�_4�f�[	G��.�IrK�����+��Y>����C[�[��zb@�â��5�4��u���觥쁗�ݟw[NO3���'b�>��P�wn��j���FƱ���}���>Uz�6i���`�H+�T���Dk r+��(߇��0?���G�۷��F�WBXcv=c�z�~j�[B�pp��#M;��g�vT�N��=ef�!�X����H�z�޺Iχ�|��E��*�UqLկk�i���Ix��dKbXb-�m)<p�U_�<Ԯ����.�)$�R���t����
w��u�}ϣ���J�~�Pfj]���I����! �."�+{ �M.�rLm%�=�B���SN���"VE�@Pk?��z��Ae��n�v���9�K9�J*ΜK�����G@�0m�{�҂��������4�"�}�Ad��le��׬	�J:�[* &�B���٠F�Pi�7UIQ�Nq�����(�UB�;c���3χ����A����q1�b=1Oy6��.�\ �i|�+F7�V
�������f R'+$Mᮟ���=�ǔ��SE �i�x�K�#���B|N<�����o�k���ˀv���`��!��	�J�&�!��z=vW*Rk��]R�I:��h{S ob@d@���~/P�w��R�`�&�a�]ϔұ����f�ENĚrĜD�J� J�SP�DL
jk�)[���i�i����`����[�!G�?���i�P���Ō ��{����)��H�ac�!Ey�lV]&b���V��_ߢ�3z?y�3�#�5��%���J�����_�c��f-G�|�LI ��+�w&����ǸGѭ�L3H�����?��ɗ���D��F��jBY��?3Ԁ�^��|ó��I�vt|J�� !��v.������[6��|h�1a���x7�9K
��7]����2ޓ�o��6e�9�  X���8���	W_Ob��Q[ڑH�hm�D�W���ёm�\����?��8p�$�&��KU�%�#���ߝ�Og|(K�/��t�/?ߛ��)$n���\��qYӁT�:G�r�$���-G�>��{q6�--X�,�8�A��@�{0ύ�n�dZ�a��O��N���Ћ�X���i��>V�$,��*�`���.+��&�LЈ�U����$hЙ7ݥ>5�cQ=cBn�����7CQ���G�b�v߁�ie�#l��f���4��VX�SMO���b$3��BB�'�
�R<�5u��2���f>��m8/�h�@q��.|���|����fY�&O�W&��`�v�m���i��I.6���J�;��(mq��r*��pɛ\E��Z��Ļ:wo�føLj�{3k��n[] ��&�A�W�HCo,�/j{�W�/Ldm�L<�7�WNqBPp��Ȱ�U.�>���ۛ�c� &�6\_�(o�C�'Ne����k�& �z��.�a�kc�x���}�(}k��9�A��M��z����~������	���z���V�JF��2���_��Nѽ��$�t� ��)m�`�/%'a���*�zi��:�u�����d���z��V*�$G�L�(y�Na#I��z��Q�BuBI'���$0����~�N��Y{�'fbGT�4}�%A��M�N�k� ���7H:���=!o/tL�!*�ņ�R܂�2���$&�9��n{��+K,�Z2tl;\�M����'�~}ɱVl�j�5�C=������1b	�m1^q��u����=�����"��4�ap}�������b��S���#���b���l��s�B�ɷ�[��_�r��	ɲ:"�F�_�:x���G���?K������:4ώ$ʈY��fy<��^�\�`�~lL�~"��2~�j~����/UH
����g\��k����}��9V�o,D�fs��m}��V�K_�c�	�m̓mʍ98�y�Fq�'r.��&����^��������mD\���1�M��z/��ݣf�_(+��cÕ�_~cݨu�:/P�݄�VjU��*�q�p��U�����2�B阳&*�u���O��ϴ�LvS�=MZuY���Pҁ_sj_�kҬ��|�b�4��hdP������a!ǋ���.z%
b�c����*Gaq,ŽHr>/K�<y8}�ѹ@���u�R��=���Y����5��3�`�9�sS,`�[�	Dv���.��ΝK��:h��A��J�-&�_x��έ��>=� Ѕ����I8x� :�`�uGRn�<s���w�^)��N�n{��n�kր^���.��K�Ke�o�}�P�����E��]f8�W���Fy(۞.�-~`�d�&E��:� <5����h_��?�������� ��?�����}�읆��{�ο��Ϟ�p>��.|���n�3�������o�<��l�FGf�Y��3�O�2�֨��b��{/n��hc������X*\GBG}��)�\����������.;����AiU���3魇C��|YS� ��2S�GҬ�X�����f�����O�EC������4W�~�ID�����Ž&�w�>��D[�j�����@1a�������t)?}嵙�W���� �#�@uKp��{������Q/P42ݖs��IC�0�sRX����C$iLF��h��	���^oن+9匼聅�1����.�mC>k�n�B��4T��Va�vtf��AƒQ���i_��s�OAkv�}_L�������-�GK�5��$$cud+����Q�;e���)`,	�|�>��,n�9˪�Igr�#�vy�a���;BX��̀��	\\�����o�,f�W��4.N�>��`�:77N��Ya�VZ�Y�F��۪�L�n���^X�=�<8��8�z����t����c���?�'���D�E�6�kv`�H�^N85��{'?� ����aW������ų�r��U��ci�<O`}͐�۸7,J5�_R#���&����v� �_e��T��s�kE��'����!��sJ�fy�Ÿ��b����6^.!�V/�(�1�t*F��M�ăH=-q��_�5Hv>��`I5��f��#wN��Uw�jQ��f7�`ЏN�kT�<��jpb�6Dt�V\t�g�z#!