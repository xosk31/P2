XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����l^��jS�wH��Ĳ���a�f�w��?	�bS���m�O���|�ґ��������uZ����0P2s!�&��%�]�{�_�zEg3�ݪG��hݫ�x����c�$s�������2m�\\�)�'�h���\f_��s�uG�u�
��Jh��>�Y"2,Ԓ焦�������hWؤ�;ك�C���j�?�3��'�����-s�z�0[�f��r���j�Ҹt����WC��A[,�?5vNh�L��1��A���3# ���E��޻���dq��Z�c��,$�&��b���8xy%�e"�4��',��-���A�*qΟ�%��?.�Vv�7��u�)F�gDL�K��G�������?���:"�����Ipi�h��je��'����U��ל,�$h~�E��M;*MrKq��h��=ڱ�5��f�g�Q���-�O���6�eRH�)@*��E��Gt*��O����-�{Ǻ�s���[C[��Kڨ�X�'�l��`k��2-�(��j2�}`�ڍ�Ӈ�aX�N�v�(������Ow�^Җ]qB�ձ��sj�w=��Lk�_���W}.�J&���'�G�&��\�b����`}?���� W�ϋ̉s15�l&��yZ��V֙,��A��O��=�sEC���nc AC��f��3t���
7ι��g۰Lz֨�:[mCrV<�5������5�]�+�&���� 1�o���w�e���|6���I&Z����'�E
���[XlxVHYEB    47e6    10b0 :u�([����47��$[�xK�i�'��R9D!+ŧ�czE�]�o�㱧�9P<�I1�D�j^��?���D�Ӷ(T`�BJ���կ�Ҷ��R�T�	��.�v'ki�>{�:�p��*�k����,G�U<���'�n��GNAe�_�U��g{�C�d,>l$���4	�����z��?n��UMMW���>��NŁ�'vK�d>�6Iք����`=%����K�;��T�)�/9I�d�P�s���[������'�S��wb~7�[�M�c5��&&zb'��?�t��V�����Ea�#;ݢ�6֣�z�=o��`ҷM5O�i�T@�v���&�$`2(�_��x������h�,Uo������%�����m�Mf�����<�L�WT9�BL�"�^X	(�B�I����ބ[��1��2���6a? rQg �o�`�6q[�������DLc��z��R��?�K�k.�-�U������)fLZ)��<3+��Ʒ^�v�Q*|VGW�N.ç��A��`��ݨ�G!e�C�p@}���eS�����՝�G��m�&�,� Y|�D��ɲ3݅$�J˞\�cEMl��e]�X؈Y�*^C��'s�6U!�U��ҨX�����S�8�`N�ֶV�J��7�M8ճ�u�J��\�h�������<�ΉE��6������/�Qf	/���'�?"��5� z��U�r��ۖ�!N�s-M���Ёw��T�j"����U��D��P���iʪw�8_#JT���mѣ�Ln��il�8���l�^�A,1fB��
�uV{O����/��u0�,U�B��A�ua��qx}sJID�3��~��6Z��|�1�����d@�G�la�	BiQ!U� �&pQN��4��ǫ���C�C�7F
_�^I�6
mӇ<�@�G�Ib�AQ4=$O3=��2�~=�/R��+�2p����GY���f� �}�_��a�������!d�	K�w;ϓ?C��p����e22Ӄ_8]�g�:�	���֕|~>�"�����\ �̨u:\	�QO�)�X��"Jgʜl�����X�Ēs�#yYƎ_Z�U�Z��aD7 ?:{�Ձ�J6��Ix��A�2�u��n����
����*����rX��4u�J�3�6�[���Gd�P�N���SK��J��A�_m:u��~M�X#q�����1l�VB1���^��;��o��7g:ޔ��-�ֱ\�6��}k�>�=���݃��]�5��������k�U �]1�sV@�A��_7p�lԟ��l]<�)�~=8��y�I�.52�Z���/��a�j�Ro�-?��)?c�����JF4&�PQd�bz�� ���y�U �Zd�։E�,G�?�6� 8��##��kl�o<�����"PB�&7��۽�(��l"Y��/y{R���g��e�!ΒVl�a�+!��Bt�%�F�Q�,�\N�q�8#�H���R"!6�λ��/oҡS���zG���8He���өܣ��^n�RPMI��Gwl=��q�/�?��lZ��V��ܙPo��(O3�C�!K�|���+��ר����X� "P�����R:V*<-�OM;�Y��ʨ�7�z�֢o�*�J�wn�0�9���8�|ʵ��Xs�����LQ����/>�E�T�� u�y�5B����VT8��P����)/k���m��1�K�ƒ���{Β�9�Np�����j��B0O�&��,�ᕁ.aYъ���M�Na�E��_�L��$��Ա�x���y�Q%c3A4uɼ!y+�9��5�9Sӈ�;m�:(����wa/����>����a�<f?Ğ��Gjl�f�� ��Z�Хe�� �a]���Dl5�V2�P<{�PJ͎���I���8{��Qѽ�y�{��;y�-x��}��u���J5�bt9���{D�"��!l�:g��Bfg���G�5ʓ}-A��8%��0a小��b�`d���b�\��~4���^�b�{z ����^��$ο��d<�Yt����zF�����h��&]���s��i����.v.�8%̂(��ĨK������.PN�Y�`r?7��1��q<f9�j�e�Dc��t�N��=�����K4�F:���-�g_Y�I�����ߚ���+[H�_�٢^������{L%��(A�g���~�Ն(�8gi_2��Y���5�v'B���FH��?#d:��\�?m2:����e Q_���aR^���\�d�5}HB�w�)����NZ���<ivؖ~�T �yY a&֙�T��1��jQ�	��}$�7�d�b���9�>)�b�i�)���i��ӫ��5F�G��1sp`23�J�-hWM�C?��y��Э�#δ�v|��v��:��NW�J�
����2?���>�|K���Pk�Iu�!��S�b�ʭ�Z�\���P͋��Z�c�΂�č�L�*��d���\Ah�<g"v��V���C'V�*T�턮�s��Y����y�n�T
�
6Q��L�nZ��Q��\�О:G*�	V>���mP&w�L�!�������Y+�V�[�S,��>_����������&i@P�!���FU��T&a��޹���:�<�����V7��S��cf��wT;<I}Yi�	$�bU�]���F�C_
��;�]�p�}�����x����S
���� A�}>�^�7�;^Q�@T;�Tt��7�
�S�q P�9��W���Qܐv��b?�7+:��%o"�kr�y1�(4RZW|q�RHH���xɎ�3�8B�Y������##��c���k�{&I���1�l�3�$Rd��D���p'���~r��ߵ6�CX�*����fI�[VC�~�l���p�����'WѼ��_`75���̞��������b4���R� /�P#rF�avl\5)Kx��`_���QR{�h�M$��=���!�"�ٵ�3ͻ7ЩEZgP?�B�{��х���Ω��z�Am��Vƶ}��	)�Q�\��b!&鿣3�N_�Lc����|�Ny�?v״]�r��!�r�a�^�"7��p�j��c'�j2���eY]uG�O	��r������Ԙ$�t:X1�`	&-�����	Zs�StɁdl-� ��WE����qe�^�K
̇�+A����J�/��Cc��%"~඀��\����������ޘ(��0D��@�J��!��,w[�]Fމ�C�sI)�S'�̶��CK`�I�����l���c5
�x�{j8�"u�Y]j'���An^�@���CM�T%� wj��O�P9����2+?��Џ-@RV?�t){G�g
U`0���i�$h�n�N�x�k?,r�����ǀqJ�B�Ys{f�:I7�,���J���{�}#��?ט#Qn�H{6�T��#y��um�du�V�'�e2�i���3(��������+B-�溜^��@W��i��h2ֲ�(@4�=��:�L_V ��Y�YX�T[�3r�5�����Q�����y�6Y�*_xK	�'[T�c�.��ר�a�U��J9�J�"4J�E��p����Rϥ��yxg�]V}�	�Ycv$Ԇ�E��-
״7����j�Z�;�������v�}@��^��g��@��K�s��Aߔȭ:�E2�S-��v��i��Q:�(�?�H�o�Ъb>G��V�ƭi��a��u�����@�a'�rP��|x1J��� #�^x}�~	tC����(�������#�����b�8��l��jq�e�'0�Z�R�}d�����HՏ�+�˖��BŹݜu�x��.�4��%� ,�rF�ۭ�� }t�$,0��g4��I��r�Ǆd�X�����n
���Ҝst��n(g5�J��i�I��yEܕ�!�?Ky��Ǻ9�sm��񬈩��2s�έ<�컢�Z�V(����5V�,�U<1)��0�^W�L�z3���"���(�0����Jp	��"�ӡlSU�z/L�v/6���>�J�5���*����^��.W�?�h54&xUN�Z�ENV�X�������`x�.B��vϫ'	�3 -MO73�j�m�pi��(���x�ߴĽ偲�ש5�k�2�aL��0o�; }�&�z�a) �B�@DOB���?�x�����y�Ⱦ���Q�3�፽�'���]���l�H�g�V�Z������!gdAI$?�6�