XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���3W�D��c�c�:zuL�l�8��YP|��V��2���T�L���xM��럔�\�����b9�!f$�"Xe��~Fn�#@:�1���q������y;����6�e�}w�$%'ܻ�WІ����������k���D����
�_�2�,��2�Φ}�y������"��7�F� �ťL<4�\���x�m5ʦ(OŋH��^h�f��i+��eV#1�f��Gc��)��!k�┞|�~��	�C�B9�Ƀ�A?xA-�9\���fU��`7Ϧ3��Ֆ47;eՠFT2�j�|�\ra��e�U�l���Z��k�^��ګ\�)b���[y��I^ ���[����7|�����y#E�t/�Ie�8�9Y�Ɋ��&]��[���<z��G���3���ځ1��gYt$[Wغq�����j��)_5ah8��Fp>G��n��!�
��K+H�u;�k��4-�~u�P�dǲ�7Hs�v'�5�����ld����Z������.���7�2o�S��Ӥ2��λ�xT�����\`x1�MU4���%�7���ʟ��b�鈁d����"�\���a8�X~(��ڰ�V��d�� ��O�Vl��zg���t�n�u#�&����XFڔ\[j6"*߫%���d&�>������{��L��(A���ݔ$A{4��_���_��w�@�h�i��q��!YI	�����#�q�+d)�1�
���U����Ų��nu��i魯k)XlxVHYEB    507a     f30�Nua��D�ə�-(���ß���B;�;�n?A�t�ǎ�C�[�h���뛢#�* 9~e���'�ygȦ�"羗��&K�c�������2;���}6G0��{��Y2),�@t���FC��k7y+f/bm�]�CUf7����ڄ��l+�K#+�i� D�A0!�3osx�N�:�6��aI�-�ۋGU�A!�^w��[W{(@|H�TBK��h��A�.X�W39�{��7=7���Vtՠ��q��Fl�D�(�8�w��L]n�F�:?�S�oo7���#׏,���K�z���e��R�W�4C���>p��[���Ƿ�C�~_6��0��^�����\�$anu�����7��v+t��Vv�-�&�1��{�hx!ȱ�D���_�� �Q�vն��D�=��!�<l��bU�&?���
��(/��5;����,�r֟UW��y�8;�x�/����{o缬���n/����4j��?��������uW�]���3i�/��nK��α�t��nH�����VKeDj�I\Ĳh��ڞ��.�Yn�69SR!uJ����t�'�,k��У���ޖ:`�r�v�j��G4&L�?Ltc����7�~�u�����X��V�R�s��jC���B�l����	��AVk�C��1�t�p�TקD�+�O���ux{������dQ[�퓇,#1QBu��	�(�F�ƶ���W6Yy9������!�bc�:o?����}Z8]���^RႠ�GE*~)��n�rP�%���:L_�:7���H��n|y��J�,!8�6��z��PyE�N���@<�gNr���@��X{���GO]
=��ɳ~nnA�ʎ,�&�/,`A�S�6wN9;�!m�����ȸ?����e/�������'��b�����vq���x8�f%; l���r@����i���?;h	iái�S��OBH���_�W�
��o����A�sg'�J����C�,���@��qQ�j�2�Oȁ�t*\n7u
�Awp]椘��0,n�C ��F��/r�\ �H�V4#�.������
#k�O��7+Q�&CzS5W��P����ꬎ3��M�5k�F���>0�������'��^NX�{�^��[���� ��r�E�	%=��A����{��VL�g'H�/*1KNaݙ���\�'�&�%�A}�N�RM������+QՆ����j�zL�~&�V�۠6�ʹ@��t$v7��� =奅b��6��A���8�~;X��Ϸ�o�ߖi�?�v��H�Y�;�[~u�Za�7J��;��`CZ}m���W���g'�=�j�3�R��L:��v~R2����Ĕ8/
��k�M�{��A`�f�-�Y�Iro�UBM����]n��1�:U�m�w[��C*ۀ����f�Q~vKv�Z���%�ij's���eY��k�M���r4��^�	�D����Q��<�C�o*�i.�=���\9�/�iʝ�'$E�i�i�+����d���%�V>��J]ȿ��=����Dy�v`˱P�pp�,,b|�"ө��u!�:�^�|8��^H�S/����lҺ���	μ199z�Ωq���뿉�~�:J�j��
��5-��,�BҌ*3�)hf�a$l��,
��	�Lo��<��uxA���1�����{fU��؄�Cc�u���;9 l��p�,¡����2:�'���A�\�Bz��W�[��cDʘ��#�G�vK�N�4�\����B��{}ß�ȅ�3:���gE4�PI"'Ɋ�&P��W���p�@ǌi�5c;�$+�=�@S����b{��=p$����Rc�9��Bsz/K/MT�.�j���*�*�Ѕ&����� ��e�ə��,ÏnH$40�8��l��N��1A����0�3I!,pu~혲KI)���j�j�ٺ3i��0^8����d7�\��I�3��ԁgV�{UV�e%���i�OM������뭚���P���v%k-A�gg�GK6-(ìۺp�,&?�Sޑ��ު��;N����~5ִ�~Y�+��U�hr�x8�RS��gB:7fWN�2	�� 6����9�_r���l�.������I]�T���!�������0�H�� p�����l����9�\��A՟��,:DQwEt�3���[M�;�Mo%߸|$A=8�����"`�DR����,Ƅ�ާ9��C��8oM�zDָWm0{]�-4�k֥�x��|��O��Z#2 *۷%;��]b��$5LPG1t�������(�Ѭ��:��:���"Nng�n`tPv4n�@Z�-�g^�E�W�տh*�#9J���5/��:O[��F�Uyd��m�>u?����./O�
���n�F�t�f�(�]�j�Ք:��~b� /����YQa��/�F��f*LI�*�[zs�t��@k�\_��,_=2��GmK(%Z��>BPj��y��,ߙ�ŉ6�H�Ǒ�o�6�A<��MM���g���s�~9QQM�ܟH�X����l��d���9 x����R�˓�2�Wjq���.C=.��Я�eC��-�F�ѱn5�T�Dҹ�������Uc_� s道�A�P�i5'�v~�Ȟ7$��"�
�n$�Q�b����,��Z5���B��i���!#��h�@��bဠ��wcC:��7q¸�-�sRŞ��5�� �Xb����
��>�jB#Ʋʺ	���,{+�/�('{�O)�i���Ƈ�j�{�M�s2,'s�~G�������JoBĜ��R��Z��5�;�M���t�}D���z�ɀʨ��S�(�s��s�����-&k;���.��<�{�-f9�J��b����5�q_ �4Y�C�s�1�\����\�I8MGzR2�]U9[��đ��+>� ?��Fe��p_�#5�ӧ�]ٖ.I��s��}9��?�_��6R����Ym�#��01�.����K��uu�@�x]~B��+�_�'S��j������?�U?_���ѰM&��E�!hB����O�Z��.�Om��^K=�+�xQT];��(-hi	,����*5��,k�S��1��L�Y��������,����feM~:/�zxOC9��B|�ʬV9M��c29�����l3$�B��������kF�NFg)p���o[�쮖[�I`�*IC�q�z������L	�����˷z?XTq��g=����W2����):S����~N�X,+���S%���?jZ��X$��'s��H�*�?X~�eT6��SP�M|���hj�_,C��-��{����~�UP�O;.S 55���X�+/��y���/vc�7aDiU�O���`C�!pWd��T,�P�֎�/���gK�2|��F�ה8��b#�?��[�Do�tE���p0Z��Ql��a����3�IG��mly�aro��u�2m�)m�Kw� eqtH�W�=�_��o^�؎,�-�T���ی��HvG��G@S(��
�N�f����3���<#gt�2�
��.V<StR2������K��.�����{\Y�YTu�{�� �^!��:�����l�����p�yS��Y�} �|���hq�z���-߰��!ؚQ�W �R��]T�	�ƭI���cz�	�f��
bK��'�sʧ��9�±X��5x�M�Z���������RA0�E��nl���G�����6��wx��?;��Ca�&}L7:�c��8l�O��7i4C�J�n�J6l��� qc��2�	�c\��L����Y!��;�3jV��#h��>C�%������%bT��m/O�q:�&�u���"��»ݺx�|�&3�e���ԟ)�{�y�&D��dx05�:�