XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��c�W�[\�S����;���BC��~�!Hj�̚�e\�II}sn"}[u�g��+B=P��RA8~!�p�<���^�y߽�7e=T#㱽���v����ʉ�mY��r�����f�Ӟ��ƹ�F>p�����g���������7�72������+��y�A���T5�2�Q�5�Q�[K,�K�.�X���-yW�#>����H�	K�ph�Ϙ����l���62�;z� �gDߺ.�1�	���� �[\��a\4�\�D�[�#�M/MD��aN�f|yZ��v
��+%&�G�r/B_`���t}#�2����+�eB[m��9���E|�.�0���7�x#]Hrs�����i0��Qa����V4�.��;w�B�Ac��P�Ǣ�Ղ-�J��[I���[���g�� ����S��/���#���d��-��8��^sv�=
��m�T&EbV]b���`�{I��M����=ق)�j��O����-
�����R�D����j%�z�%Yǹ�V
q��ޅzY41 ��H��>���(ȱ�4츚��NI�e D Rw��vz]0,�?�ܘ�K��X�c���b[̓�����r�7lVC1KJ��L����	A�ξ�gW�Mҭ$~��s/���1�w�e\t���Ŷk�a]���!�jRH��lK<�{,��[�1�[�T'&���YT��A�v��N�D���jY�P�B�tX�@���C8����StM�T�S�$T.�0��@x.��,XlxVHYEB    33cc     da0�Մ�ZFh���!�Y�#g���X�8���%���n]���}����w�`�(bi+����p
'�hRZ0��Y"�gkJ!ٸǍ�i]v��㷘W�'k��̀�6w���Խ3_���ryiQ���k�ڎ�/3�B�W�H���$zm����q�MY���c�~�tw(p <�k��CЗ	9�O��U�C}����#��b�g�b�fj���>e����}D?�sx�K�a���Unj�M�A`����{D��x��zw6˷�QVV��w�`ɋ�w�$C-�[�A�֬�L��tM�u0n�q_O� ����N�����Lb�Q�2]\����31W{/���;S���=�$��|�	';�;#�A���u��^[!��#iy�e%5�/�B��n�`h��M����M]"�M/n��(-y�&����F�ʸ	���	�U��5�X�?x�*7���U���ۃ�/Nz�iؗg�7Ȱ��N`B���_ӽG���39�iz�YTS��Q�k�ҸwS���`��v#=�9��?���$��>�����B��A���Z7H�aqY?���߮-�XB��x��m�7+5ʥ��w�}���9�}�ދ���T��~7�����|1q92�ʜ��2B4���L^��hC�:�~��g�QB+�3����U��B2"�d�ij���j��I��l��]@�.
�!{�����]��mC,(k�s��j���}����x��5^70.�Jo`���l�4{XNH�6<���%Z_߈���i�g�i`˃�<�m����8L���������j��DQL��
<a�4�vt�u�tZ��g�Grpy��ٓj↔B	�-D�g���Ʋ�a٣���#�1J8=���|u�K4����� ��aG����F�4�I��vt$$L��x�̫W�1�Z�n��dku��Zr�_?�����/\�f����e>*åQ�ʘ�`2/�Ҟcl(���5���ӁW�QN&� �m6"\�H\U�͇�'��F��^5Kh|tsviXQ�&>!<0CoP$�|r�U����}�%t�j֌+]J�?(F%�e��6K�8�;��C�
_
d��,.�o�x*Pvo�R���c[:�X��hk"]�M��	c�5|^2�/�@k�IN�l	q�V)����w���Fe2�}�W�K����g�C���xh�/s��� ��WI�3h՟�gؠ���,�;C�Ǚ��{u�|��̴"O�8�3	����!�l;�{�Gw��òC�؛Љ��6��ː�����>߅���� �X&��VT�v��<�@���p�� ���|��x�W���[i�ؤ�}�74����X�na����/��l�9��R����-ch�]{v�L4v�=���BB�ݫ��ԓ�����`p?�:>@ϝ�0�����oѝD���4cW}VI<7���z�����ڶҶ�Xs�gf��Q��|��{����J���I0O�F��3)�W���C]���B��z�o�;������Kxգ��?n�������-����I@h%}%�'����� $���6�*��7�*Fz:��u�w�����W�B0����̴���XnK�a鯠&�Zy  ���<E��Pt�`�$ ��\��I��*�n�^]��#H�Q�cםո<b:��v]��dt��F���\A`�B]���vs0�CtӉ��)ʃpy!� �G�8|�dm2dtHՅ��A�Q��'_I�8��Jx�VvQ�P�JlHC'ٲ�+�ŗ?)(h�	���U^	�f?b�<Q�0_���
֜�	�=�h��;�'��RY�Jw�#�7�Me��Eƺ�f���3k��; �����"���=:���S=��F<9��� .j 53配9�����Ffӟ��&�/ mB(�����{�Y��ѾCe:O��4�x�^�Ն:KL��z��-!(�ER,,d�<���ƪ�$a0z:�u�=���_�~����9����U��Lq��e���1*񛔂.�懙�宵�|4��H
��&�Շ��_�\Y!��4�6�0�-�h���}��`o~B���<O������*J������$i�}���T��8�
�Ǒ�`�6�_���V�seb yg���r��,���3h�n^WMF[Ru��U�[�	�Sgf���\��[�3�D]�Y�ĭ�Y٘�����JM	kC��}�
(ݕQW�w/����e5L"�&���?V�������-�g��j8HWȳN�el�f�ꎰ#��B��Z�-;ͮk�#_(8O��7G� �~?DäVv~ƪ� ���s��38������K��m����)n;�
�;�PL�liG��|:��9[��y�*�����V ����,�.ٕ/��H/�;�chs:(J7 �oM{;�MjSQ���!,�0�"=}�O�6�H�l^���}�>r'
PS7������%���(�%�O�D?	�5V��:��g�I,�qjMG��Z��\��Ǐq�9GK0f4�Ai]���N�6]|u�Y��6�Bv`����~��0l�&��5�ӝ��\��!+�F�$3k�.� "�"����&��a�Qqј���+P	k��_YQ�c�?�)%�7T}�Z*���$G���&�#k�Xݑ��m��@�RF5"ף6=��g!�m���-Z�}��@��E<._���#O{@J'��,!ե�0Or���E�B��qD�LΧv�ʮ�N*�����\�q��lp�l�9��i����7s4���g�>����p|�q�'1DН=j�z_p��K%�"C�z	}��zh�k���VyEG.�����s��#�I�Ž��G��z5=To'���h5w��'R�ר�	m�A��S��k��^Xh�z\����B��҇�s�c����l��E�ݐ;y����;�O��f��N�,P�lA^*�� ��U���/�͔�,j�6	A٫�CU�����b�ظ��&d&w:��y���l\8���63���"~pR���k�L������Z��A*�HKK�1j�L��x����2��2�M���]Gޘ�ڵk2[��i������c~~��
�]f�v�G���yb7Tt�� �J·P&be?���*�k����5�O���r�Uk� ��GSݙ5���N*SF�MY$,�}k�07ͮ��w9�����z݈��*j� mn���(�H�9�,u�ǩ+��g�=-�� �=NF �g'E���p��i00��_����� VPs����}�JOF5���x���^q���+-�+G�֜�.��o��7Ciֽ�z�*�6�K�&����;&�L�ydwI��������J�3���~r�HoT�ok'�%�l<?\7�'�)��6�]*�%�1r�D���\U�/e��a}\� ����o�'xp0�\��"۳�B�yÛ2�{A��wEѯY�����]K��kE�'3���85
��o���`^n]��~��T6��*�