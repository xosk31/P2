XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��o�)�_b�C��1��<��g�9�?O����JU��� U\��M]��e�I\��V�.�pƇ�Py���J\A��C�P��3��$�x`lu8}3Z-?�DA�7�9��Ú��/ta\jnp�em��jx��.9N�O;��h" Df��l"~�Ɋrو<"�R�ƴ�����}����[�~��
$����hy<:꼉�	G+�sŹ��d����4-���M0P��ܖ����w��c0Or�\��H?�<���cUZ�z��Vw����Μ�xoQ�1�%x2O�_�Ƴ��u���Pe�8�=������:�$��F���������7������ԩ=4SW��+\!��`۾pO��&K�X��Mʁ �@����wwGj� �;���I|HN0fC3�(	c�H��m��x�<YLr:tRc��֐4sr���_n�l%k���=�>�{��g�(��P�^�
Q=�z�=�/���h���N�^�l�Y*�%�*�i�qصI�N�yͽ�Q�f*�%�W��P���- p�L�!�~�$TSzB�����ආ���W�>JIj�1Ը��vɀ�����<e��`UV�yy3�?&�q-^�z���	�W�x`���Zf�Mؐ{�$R�a��Y~�۫%��;���Y�:.��R�ݎ1���Y�ђ��c|��'��%@�r�������k���+iJl��8��?N5[D�(�{G�{�!%jY���6��؄��8_�6�n�cݥ���IZ�մd��'�Y���XlxVHYEB    fa00    2240̊��V(���ܓqjO�I%�S��D��T��
�C��}\f4�w�pt���P�/��u�Dg�g��8޾��b�8@�4�F���E��8Ub|�̇����dUn3�-Rvl T9�f�=ϺOO���}�!@�k���EHڈ����w��M��42������`��:��e�I(����&uZ����$��������I`ϧ����2�Z��vs��E �����[i/��cF��&%i�uUmV���;��5���qÓ1g��Gox�>G�j��v��͟��Os���zޯI�-�^t�<�\����yC-��@��l0�R�������k��ˬ�1�&�/~A���lj�6ت��^�4ś�42��`c��szaf�Fo���/�=���W/�i67�|pn%�R��	�5�!�旐1��_��?�*������#�z�ǭ�^Fm���^ɹ��L'� h!N� ��;�H`��x0�<Jf�+�����0h�yӒ�q>R��$1�/N�^Rc��р��u:J�NE�!�_ovX�T���[� qRь3}+D���d�3�I�˗�a��ܾ�����e����yjn�Ps��!��G!T�s�$�G?�k*i9��ňC�Z7�>Wj�-�S ����}@�ŜV����{N�>`��)�[��Y^`�i��R4�|s�P���X3���8��t���0���3��D�mh�\�`����i�lꉮkI� �NV�0U�m�$%� ���qB�oQ���.����`u%�qVzu	�?�9��~�f�f)8�V�ٸ@��RJ��"�9����%rk3�:�Ye %8�R%z��������wj��>�~<o7�����g�Cm�a��<jpN[i(�/���ׅ�������'��&-Y�7��:x7�5jZ[�J�\��?�4\�I��S�>W	�X%�=�.=M��q�O�~�Y9��L�cT���l��c�9���D�˾Fp���O���m�}�C��{ȗL���n$Z���S!�aV�|�JWDƷ�����B�����`	R��R�7X��}V6(�I2!�� ��FP��&�<O�F2�)��?�_X�mߋ���z��Z�jO|K���GO�L�C��ܸ���X��Ӊ-x�y|����b~Y��Mr�ϑ���0����,����y�Ҏ�O���}X�J�|�u|z��:h9G5ɉ���Lf��t�ImmI'\x9��y|���a��1:�U�
�r��YV���ok�Ь�ݨ�$��nx�-K'p,R:vBչ�zN���'��
�v��t���&�����S�6�����АܼYy�o*�H��
��Hw��SU���׾g�I鈳��:�@�,J��ϒ�3#���I~m�Cѡ18����] B�˃ƃ�)1�~�$����3	[�3o�qΤ�����)5J�z��^f?�	@��uY)�.�i�U�Duf5xȑo�$��B�e�I��q.&|��01����
���4�:�h�M��E�'Q�a��!28Y8;g�9���$A�e�Q!�`���S�]��3-��'�\��aIR��FXWw0�6�b/�������sĚv�9G� .�^��8��w"���\�i�18��~[\�H���4��S4/����ź�؟לD	P���F�Aʘ�8q�c�Bhbt�A��
�M�V{�j�刟�F�y�yP�w���]�S��u�쨢ݧC4sE;~��蜓�6����${:͜�g~$�����@��J��v�H�q�G��Y���`��]H:�^;jƳ'ą~��Ex�r}#�x�JX�v�����)�d��MX��W�����E�\w<��|ʑ7}�1�Hm��	��`sj-��w�Ƃ��fk�9,\�W:�z`ٹp�v����h6k*hd��-A�L�/�}!}2h�vK�Ir�m,]ۯ�{dCyfR��x0��'6$���&X��,��GWb�N|���U�OܞF�]�ᇵL[Q=���|�i��Z�Yd���뱜in�`a�R�?<�gC$].!5�4R�&�e�r�6E�m�͵�L�Һ�> .��H�(	��e���py����[ྎ]�������/��	e׶�
@b��M֕% �f�ę*�{J��K�kлʖT@w<h�_X6�`����\��ϵT�?n ���A�
�_�{ �Zrـ�rj�o��nf�����c@Tù2���j��I
9��C^̓�*�y���a�O��7�Dǎ�o���|G"�~�hx~�9$R�'��Tp{C̴p�c��I�ЈW3� (*d�h3&1�D��ޱxP���s�u�$�p}��ūw�9��+�G�Y�oJ����� �>+I�N�Ym��YO}�n����h��� xLK)���*\�̂�'(Dg L�����{o�QFme�-�P�89#�����.�,\�x���JЍ��ŭ�0g0a�Yx�т֊�엷�"��������|re��-R�6dS;Պ�]�o�Y)�Zq�X�^����&��؍���� �R�eC2e\&:n���%l�C6�ŸdyKh.��Vd��Y���߉	v�*-[TT(�r�']i�_���j}�V�/�z��,11�yYo[w�����/i`�\��#�N�����t"~��,���h�C�`w���c(��}8l-�r���3s2vH���
4>�Ӣ�kf�u�A�/ɱ�}�pi ��U��3��?��aPT�����j
#j�A�b@�-g��5��+x�_�*�v*��{�=^�g�ߨ ��*�7#�Q��ps0*)�+�������.I)&+{��Lk٪��7��66	�w�>U�פ��?�4Z�0u�Խ� �NN��=и�:��τ*K��Kq?߿7�}�}�]e��<jo4�~Q��_߄w��;�aїl7%cq��#����m�aL�^H0��?�=�b�v�<.��� ��q\����X�Pn�x>4��ZXC�@%�Ւ@�C�1_*�}�g��tw(�����}��rJѤ�q;��Vi)����`���� t�Y�W�㳤�E�t���;�3����AQd�f'�S�l��^텚�Ex���ɭ3ߠM����ոx̫�W�g�V��{$>H��R��%ve�=�C�cu�\��@�
QoԮ"��������v=�NDFa6��9��Wl����-���ݚ�O�G'3�y���I�@�I8US^��}��y���f�njn��o�{�뺚Iu��	���z'D�1H	�#_��.�j�l���ګe����Ɔ����X�]�X��q9FC���<���`�s�I#N�)x���5h���(k��%F�l�d�DOZ�g%�Ky��2��s��1ҭ���=n�""��n|WT����]|�C���ań���a�ԅoH�����+j��3�U�O��<�AE�b�L����=��W�P��Yz"k�˫۝�uq4Ƣ��=��߂�qeۨ��(m��UO���=(��8 �H����B�N��W�{w�Cq�Q�����^`�w6�-jceK\�`�8N��"�DS�i2"a�=WV��:(L�@�Xߓq���E��j�MJi9�)�,�9eB��4Ms���e�2��W��>�����ߡ(Pm���m���.m��;�'��I_�GM�<��J]�T޻��#�r����``7c�9S�X��]%�*\�2^���� a���b��~���z��$���w�H6��'���/pc��
��Z�^��Ĉ�_���l��Q�)�J�G�>��MN�Yl���ފ`Dn���c� @h�ӆX["/lUӁҏbЋ5P�<�.r��zH�,ta�J��k%'
}E��	�� ��_<�h(
o��8I-�vZÛi���]�������4`���>�ޔ�)~�*�B�Kː��e��ѥ�T0����.�z7�C���D}/j+��ߨ�gE�|�ez�S6�ұB���f�%��=���͆`:�<�*���h��=�A�rב�i����B{U��P��׿�^�)�],�XM@jL=�l��].��E��߳�hܜV�@�cƤ�%x�sR�h�P8R���f9v�Y�	Г,��H#ִ�E�Q���dZ��87����??O���u��%00jnܒTg�i�3܊����Ru���&t����"��d��,2�t�q��|�-�h�K����)Zc'ٵ]�T�4��\/���-x\h^p��5�P��Ev��甹ߍW	�[(ˑT�=��q���/'[���2��P�ڲ�Yw�p���\��:�������!�P|��=0g���R�>S�Y8�� ��C Q�ֻs�q�$�ް+���}ݡ](U�5S�%*)��O#r��gNXy)�?C�e]T
Ԡ�����R�J��ݕJ�����.�4�B�VU�{��>B�?�� ��<
��d���Ž6�Y�B�#&�?k��LCI<FӢN�0����Uш�&5��OVjy!Vx(k�҆��8[ ��u6� �l��`�D�@o�j�\�@�|���V'�c;�c��)��(	X_���et� ���"I�Z�K�Q����4 �p�(�+$���ʣ�����N�CUN�w2�ti$Ʈ��oj�u��z9Cïho����EG����f/��?�b��T�P���L���k����6�G糮3�<��\�	�,�Z�}�0��E�9�v{̗�ֆ�ҧ=j�����3k�ԙɧc]T�bA�d?�i\��K�ջ��;pe}W���2����9�tN�c�B��c�3e���zoM"5i43�C�1Lea�6_���(���g(X8����1{�tt!�h�ؗ�(��Җ��A{e:�lV�z������d0)��egϪPA>�>��\�O�C�gk�k���2zB���%QB"c�]:؛��C
�,E�=W2찰`�ͩ����R�b1)�GA��æ�v�l�[���|!'Wk7�g��w��a�F)��&=SK�`�VD����.��ȷ��خH7��_eE`���d~F5��B� 	�ۆ21��\ƓG#RJ�o��mz�
�o�?^��D�l�`PV�H~B|�m'�}����埝.%�vH i��/���Q4�W�.��o*�NL⻻.y�Ez�SV]�Xљ՛x��!�e�2aCb��8o1�6\t]8n�.��Z��n������}�ҳ)'L�'�������8��U���<���͏�٪)�cC�`í�X�<��æ�9�J��J�g��"ʼ�|��/��T,d���}Nm4*񋗓g0��>-��D��DG��o���:�!�(��Ԯ:/C�7Ak�D$c\�ܛx��@����5�
��/�����9�8�.�lzxs"6T���f-]I��T�=��=�7��xB���^zh`2o[�|^Ƣ݇�֡��8���s��U��;�n��a7?!��Ɂ]��B�v�dS���90V�r�&	j��Ӷ�<��Ts��Ft=B5�ЪI�_^}�q|�9�T1[���Or�>������xj lo�A�q}4�4�Q6�\���%gl�C(�f'��=e!Q��TC���z�$u�
T�t{Ts��� w#�)u���L��PT����Z)��k�9�X�Q�G���՛�s�Y/V?j�����+R%\^�쉷Hl��襦���'��6�F4���Z�cW*^��r�m��YCv�{�u�GO�j|�@W��ӭ��z6�:�.�}�iֽO}#�E�s���4��A�d����a�����k��w=�4Y��r:���0�⎾�]��[
���Ӄe�&�"�BaA�A[�iϤ��6�P��Z�{��n�0�zbA�g��]�k�׬EB�L��c�~>N�89�N���zs�GO��!�N���H��	wF!�'���8_�G5I�������O�f�����F�v����Q<��F��/�f
Cڂ=��Vr RR����ՠ����}��t���jh�s�yO����X�D5y̟�W eCG���a����b�̦�|�l�޲n�`�]VwAì��=���������R��-�y1w=���	���YK�Q�/+��
� $��鳴��P*v.�_�C��8�C��� UW�Fjed����9P���%�{%�X}�������0��][�����?6f�Qw�q� &w���;�C�QX_�Y1D�q�)H`u.����bd;�)�C� ��!!�>���P�e���};��_�bY\���/�: �s��_ӝUn�юpV��$��#�o��u�.�%�.[{�>t����+��Hh����_[]�e�n�-!��aU�ݣIv����c:A9�+[���� ���,^qk�a��&�縛���E̢��9���8�q�;$�IMMW~�}/|�㌜5���M~��/�B�;U����J���A +�p�/�������F�fҞ��  ОHY�MZʳA�sn0_�+�N:hC̉]
���D�ms,#
Q�i8���g�b;�[��n�a�藧��O�E�Z�����/|	mH��$�v��� �h2ckP��)Su9=�?ϖ�%�F��$D\�OZ�~���KF��z�Ƶ��h�"�k����"6P+�r'6P4ˇ·ӷqV���L�%;\ޑ��S�QZ?~D��P/���h����}!��p���D��	q��A���Ur�-W�Z
`i%�K���'��_j������7]�T[Iuf��+������0�۪�M���qR>�9;D��Yr=+�u�9]��7`6,O���)x���Z:���H6��)\��_�s�zwc������-�����
�m�����gZ0�2)��G�����Ҷ/��O���	}+%�@#���EY%!I�9w���FX��g��f�m��t���y,~�$�E�b}��_F������Z���:���twʱ8&h`��]�
vtO���[�*�lE
%�"~q �!�0�v-I)�ͣCv/e�-�,����#Q���������!�Ѳ�&	F�ㆣ�z1.�lMs�;��cZ//�@$$��_��Ѳ�*i�s�����?h���޻� ���9��b�W=�L���+"�i�O��)��k���g�F�c"+y�5��M�rT�K7��}�!y�S�]5�P�G�	��xߝ�P�@S>J�|�{����Bn"Uo1�����8�*�P��2���r�ҳ<�7&�#Į���h�f*���Uߐ` ?��~N��@���~m��N�ԣ�"kF=�qYx[-'9�����;�Ux6�M�𵂺��qk�P��� �/���=�l�ߢI��L�t r��3�	?�!��!Ch{-���>;���e����I�e������&d���l�&ߑ����J�	���s�֚f�g��失XW����UJ���S���]���>�V����܁?�`ޮ+�u��d���8A�Oɠѫ��ڢ1�?eί�G�k�.+t4K��Ln�À�+��aQ⎒�f~B��z8��rt`g�֏�E%ɽ�)B*g�1C^�i��$�NY��F��>�V4���;�O�iK��I>"LN�(v�|��>N��9���Kj�@�H��K��|y��`d�y̗)�H)QX�d�|��M�ۉ�{�ğ����g��r+���[yQ����U �����v�opuR{�(~M�S�\�nʙ�{����DŻ+�hCN߱��*��6	V0+թ�&��ઃ��\��*O�3�����+\�_A%^I4`4$:ls��:��X(�|i��rB;�X�+E���X�BD4��� �ş_^:d��ѵZ���R��+��#3g�{K��M���<U����2D<�ri��*��s������̫�PCt���io����
 ���U&{/�ˍD�d'�_�_�d%���ht�.ʬ��I����75B[0:.�꨾����`Y�%�^�mɲ�����!Љq��L�JW����1�eap�NA-��h��M�-gЅ8�9�����M��U��Q�+ˍ>��@�̒	Tn� ��'l�&�F5t8U�~�R�q�wScQ�l@���w7R�����k/�r4v��a���������ưNHk#����o���w���~L=�Ե/<t:	M�)��"��,w�/� �C�c��3'�A���`�l��:�1ۓ����}�5>���HH7̗|�� $��#E-��u�n�["
�	R�a������䇣��L/B��l�"J8�.�CZ��Ȓ����i�
�f�R������WΝd��#�ڨ*J~)dp߄.Nr�53P�g��c>�Ku7�α�Eͮ�����ж�pbP���Ŕ�e��wS�SZK2D<f��"�YO�Ru��E��W�쑈���a���{�뻕x�t�(<�w���9 � [��qjv�SE�kk]n���X�����΂>�*+�dZ+%>4S؆f��g��(:l����݇yR�$�5."�*l�|4���܈�G;a�v����wq1T;%����LK���6�����J�0�ؿ�G��O-E�w(���L�WC1@�$j��^��!|�r"SV��}}� ���{`K�j�^w��L��x��a� Us�^�Xئ  �t��TqYw�>x��!��<,BG�qv�+KE�*��ad>�Ӛ�*�60񷾡1�t��@{�<����~G� ������쪆XlxVHYEB    6682     5d0��5qo����a�r0�FC` ke�Ҋ{��!�.I q�;��'��.�1�le�xz۽��?�")jEa��2�����>�Mː[f�z T��M�Ȯh:�Ԇ��0�[7\�������+̈́	��S�h�BY��O I�&��V'I��_�����J�����B�(��M�i�U��%.Ћ_dg��ltb�׃�gwY�a7����~����y�������I�_�A��ns6ӏ؜�yD<6�)����W���ݴҡ�b������A���D�0�����Gw����Q|s�B��&�&�y�=���(�j�bv�>����>r�mG�%�Gk�H���T	SnT}˂�Ԍ��7�E�U����s2���0κ��X����;�_�G��4��!�GAL�j�m�J4��l��a@�7�i���S�+Z}zf��֛f/�uG%��.�Ĭ����0d�a�*���c���R��w���:�.�̕�-�J��fAT�M����)�+���B��G�R)�1��T��� �R��aCf�`�p�����23Z� ��)x`�;t���	��#�_?�'�潛�!X�j�O��ip ǻ�#b�D�_���.�hp���H3�f>畈"%��2����'b�Ʈ�Qx┑�.�6�֌�1���"�zŋ�xn[{��:өtA��W@����`
Lg�v����j�x��])�N��z���ݥ1���>��t�+;Y�J5�<q/Jf5&]SM��'�e�	O���S��S�n�s�{�V�	���5���ΧTeQ�e�S�0������K�L��(a�@�嗈�|	ZC�5���q��'DߞԳ(+�P�C��z�������?�m� Q�}a��}��$R1܀Z�8[�s���4����j5`�u�I�,���^�/ufԥo�릨����S4���z��.���/zTT�T	�d $;������+�!��h��荿��8�5e���P��%�@�\�kd:��X����p��p�6+6���"�a��Nt���(�� ��&�%�(ĝ8h����K�g����Ǻ���aGõ�&.��6τ����d0<2���n�&��ݟ�Z����1՝��<a4�5`o��Q3�ĥ����i���C��r>�Ϯb��P���f��ԅ6��ue��Z����a?n��2�h�����<����l�<�n�6��bi��n��J� 
g��,�#LU�i�0��0�i�$ܯ_('ư��I���F�b�ە��_��vt������yh*^���q��0�8��Pf�����}�*�֢j�$���$���)��n �dn�ܭY�.zs��%W�c\�%�0LE����ڌ�(�!��D�]���d�&��ca6�"�x�R�������;ߝE�>jX��_s�zy@ ��\�``-�w7���,]\<�)�x��q{�l��x)��C