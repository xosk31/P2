XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��{���[����f�p��q�T&<-�ZC��w0y`�WHt����p��Hq��3� q�T�)[��!V^_-���w�!�p�e������1����A�@|�C�6��Cv�0���JP�d�*�kƝKvY�,O���[�R>��r~9R��](>�].��a�����2��z�)Vwxc�e��Jr���Ό��������'L�˓�"뺆ϑ��TL���=�,(�� :�p���2��:a�=��iUp�A�~�n�J����J$qٖ�+b+�{�M�K`�V|��,	~���@�kZ�����]+�+�����>�Wr�=��=�l�7N�8��,����P�Y-os�y���0@�]f���]�.��;fk������U&�W���/�-^�]?�4=$��m�v{�_�m�|3E+x�� u N>(�SOZ����\[�,3�\qW��8Jym�e~g���aU˞A�K`H��b��8�U�� �L�@��Q�Js <���='q��w�A�
���D�`�M�����V"��N0Ѻҟphm�N��/֊z�N��sP��g������X���YJ���s�W�jo�!C�4P��;�T�]	L�-�?P�%mm/���$�� �A�Xam�OH�o��1�N�qs�`o��1���N���qf�%�4��tT�LJ��u-����y��:\ �� W�u�n[���
d8Z��P��'��TUmg�nh��ͫ42"���;����l���Y�y���W-�
#��8w�n�+<�ot]ܪeXlxVHYEB    9efe    1be0[w�#��ayx��M�8��l��9���&���?2G��!h�M\�bMy��@����-=p1KH�<3�3�a�,۬D|{���5���u$��f�c�$Cʰ��i!��H��%�3vG�tanZ=�	��|U��lWG��h�u�ƍy��\�[�P5E��*� ]ƒ瑞K�Ҳ%��؟�����,�Nk�q#cuiA�
��Q�h�U����(�۽ M�w���;�k	3ܺ��m)T�0��֍E��-fmU<Z lPŜf����/J��[��č�,�b7ԋ�#��}qNL�.�&jT�1�3J��:��n�"��e\�,[��l�d�o���*t̐߱Y��gǦx^&9��'���ݗt�L�	�i�i��;W'�څ(��(᜶Q?�4��~B��m�h�8Y�# ������!zc�$~0��\�/+4G�A9�	t�ɞ���H��4h-g�ܕ���R��0��~c����6e�Ը_	"+����~Y8���A!h�bkG1��]΅����L��(+M/U[	+����6g�D�6�iH�6��	�`�;ՐV�@%��\�v�]�5ĺ@D>����V"k�+sBgH�3��;e��J ~����BR�ͳ��RY�^^����ڧ�b���c���hj��u�f9�&Y��%+��+��ER<����j �����;�[v��N�iM��"�}$[7�L��*�3V�6��t�U�����OL��
�� ����Zj���~\핸ß�����6��<M�2X�1,�
���Z{A�;��6.��b8\���j5�$A�5E�%�	#��jX��*�MCF�(3�?@��8?,B�t��d�u��[=ο�k�lQ�M�*�}g�xN^~��_�b�|<��ȿӪ.�i�S������B�{�7p&Vo����%S`M��S!�� ���:3T�".���t��)��P�О�TP#�`�zRW6�ϙ�Q�8���I���?�GW5L��px��a=�%k�Z�~)N�e>�J�&���2�7���n�E������̖�{mV�������]����dh��m��ލBS�l�s������;�Z��J+;4�XfX��@+�S�8�u�'Ѷ@�d�� duր�%�Jj8��c-�n���~�AУj���%�ο����n���U d8���or��܎,������IÏ ��S�O?m��{C|��y"l�M�\.p_\#�z4����IN*���y��S���,ZWZ Gd�A(bd����Xޔ�X|�A�=�0�(U�#*�KG��&�Qś�J�~'��	���܊�5f�"�8�i1jK�����!�Gr�*0�J��8�aC.'���锤g�Z�n[D�e[��d�
�?,���nE�ž��;qe�c)AIێd�8�3�;=̂H��.�.j�d�8H�_��p��}���ܷ5����R�hEw\1s����ч�p@ݞ�Kĝ�ܓ�1vh '�3��G��ь�����=�=�yX�ք��1��5�o�"��������l�) RP���B�}`�Jh'q>Z5�\�?y����R�jY�!�E$b�!B�O�8`\�@�ܭ.l,�Y���]a����{y��7-u���P_O�����1�M�����cs-��/1ȝ|g!}m���ˈ���+ߦ[���ξc�s�f���G3M`}8�k$�L�9Y4`a3�eY�dmFZ��v٣U��+�G
j�sG�W攬�J_�C���g�j��K�'4��Tנ�-(Վ�Zf�+���/�����Q��>�YH{E�zV��Z疛N[��l���2��D3]�&�!�7�9��ئ��?��N1�s��/��oHB��p&�m��_�|[���N����C%p�4�٪a`�ڣ2����OW*���ִ�6��괵��Hɘ���1R��`}&:������1��ȩ��D ˅q�v�1z�-����a��e�{�g�Ru@�c�dl�:�L��ױ�[Q<k�x��z�Vۮ����J��{U�Z���S�����L��"�Е V�,��i1rH����[�@{9���ۏH�~�r�؍� �����6����������'ҐyiK��IG��0'2�y���� �Hb���b�#g����u�#�O�#%g�?�v�%�qL��� I�ԍ�YAieT�������-������"lk�M�x�ͻ����F��`y.���(^��<�+96ch;v����nX/�����p0_�ё�Gt`�y�X=�٪���UN��P�� ��;�k�t�K@	�.�&v�#�ib1^P���Q�Q��Ǳ	�'�� �]o���H�R�n��%�6-�N$P�=y�WN�o{�%d�B�vg�m��,C����j�GcIh��K��HR"Xg�QV�\;[��0��pi"�l߷�Բ�G ;~���Zb�VN1�p��>T�.��G��x������Ҹ����\��\ۖ��}a�3Z��]�n
 @�5�Q$@}�-�B�s�50�e�#V?"����w`63L�=�d
��L���i�5{Ι<�~��[a����;��X�'�n5B��K�Q`>���{�2��ф���R�a��*�O�Lm�����X�1��c��ȟ����t�@�1^�<2��[����;E׈�RR2H��)γM�43����+Ȫ=7F[���\�߃���q.	�=Q4������JErm�=H��M߁J����o����W��C���{�>�<�BS�g�v<!��W`mtRU��������2Z��s��c�����
Tք�ݥ0�e��?yhצ�á�҄�b9�a�Ι��˕�/������J��&Wӣ��/}{����Q�`#'[F%3�� ��$�Z��΀X���e�͑<:`��{!����.�7,�V��v�^���D����5�*�l靐�yܡ�*Ħ��;�:J(�e�^=o��#,�9ְ:��Cd�v<D+1�ZE�aXPNi���������g6DDO��^
�^E���|�����m�QU��f* eu��L�f���k�i2)c�	��Y�?�׍v<�R,=�=�S���-_���V�q�3"_�_��q)Mǵ��iX�a��+�h��r��4twf�9Y��T��bWe*saQ����:l�8�`�����/�7�/�t��DKڨ���l��y[�	�/ArI(�a�p
��<��H�1y�X�u�oc^�f�|B�&ԁu��l��pS��<X�G��D�ivb�����^\ �6���]]�U/!�r����D� T���w�p������MO=A�g?8|�-�zJ�2�$ծ�Hr�$./�>2N*bT9�X%�hI�9�M�OTL��U�j��ѣ�6��<{&X�z� ��V�o �D�[ށB�VѰ����r�x7����[�B�+|���	�)�����]�S&0gi���3#�ˠ`�WD!�J?�s �,"���&�����_�hØ��ݰHI���Wԏ��m����/���q$�O� U�3�����zb;�+b
�q!���1ԋ�`; !g���^�����E�����Í|���r�6�R��tï�l��/��N���i��t_#�,���{S��-�J[�э��cb��-�T��7�^�5�5GթA:�T�l0O��$����y���GC��>7c����U��2�f�y����|���-U� ���+���CTѸ�UK֡���� T4S��(ˣ^��A�IZl/0�3�h�PY.�D[֨$o���H��^��ա���a) #�_g�FUy��A��S8�G�>f�t-��Z�]��8Fݲ@���+�*��Bp�u�eܻZW=6I��8cLe9���� J�}Ѱ�����	/�+���R��L+�Pp��rt�(�!�^m��r���zܤý(#Iˇz�o0ΰ�G���|=����đH���δ���ȑǸ?��2�mx�V��L����h"�����c���CI[�d;��
�yǡ{Awi�:�!.�y���l��?�ƣ^{�y\B�m�۾�����YmQĦM������Mv��w�3�u�8�Me��1����
3�{������Ӎ��<q�#�3�gU[o��I.?ǯ�m���Cj�FX�7V]oѬ��+q�^F�	g:���6h=�"��&|�����$cUGr/���v���_�9���J���!���`c,
_TK�Nt�ν�p4�\̨���ͺN�S~�Tߔn؍�+�6�}�i<����*"z����3C��<8M&/�n{˕���|:/'�d�T���R�w�$��K<��?(���W����+J������H��gƥ�q��:�"�w��SR6ʶ=��rf��q/�Lm��=���h����Be���4&�:"\�N��혪�-
���ja<�C�2O�w!����Nu%�a���>�v��>�9M�q!QV�-��������:k��"e����94BpB�������9��q��i��Mx>]�ޒ�z��+��>���r[}�����O����j��U�7�FG�WQ�D�,����c�:<����賬 ��Y�A��[�>�L�O�2̐����.�cn�C��u��KA�X$Љ��&)@�#;8�f���Y,>yƱH��0~e��T��}������|���VQ�PCpy����io��; ò���?X�T/ ��Z� �*�~�dA 1�Yʥ��ަ��rU��*p�ѝ��d^���.ܒ1,��9�Q ��3�k��,���#ۼ9�M�x�:b�ՙ�FO���h@�C���Л����<-?�a�s��Mʚ��ޖ�k�{��<��G�C�6�pHì��lݜ
H�ǿ�ֲ�0��N�lc'(�3�Ls�n`�wd�
��+`J��%M�<П����%%V}>�Q���X[E�y�Yw껖��R��V,�]$̶B�Hyϖ��ڠx�y�d�������}!M����[��"0c��ɾ�Yo�ˤ�5G!�W�!S��T�F�}~鮚[?��������[vɒ$��M�A�!�yH\�à�~��5�>���j�ې�DY����X���p�����Y���>���$��ѱ���.帏`��W����s�?=Mj3��w���j���c���N��5���X�(�<���V��y�Qq��vx������rh������o8\�&�jyd�z�+�d�	P���y��Cg���(�	ί�C�ϊ��Tv�����s��Ɋ%K�K˄�Q��.�=0��"M(�V����a��p���sF���~����+d�����4,Kv�b?�Bd�ޅs�4��7��2^�Inш3�����4�v4F�	W������2(���r0��e5�W��r@��~��ZS����f�өϟ�)�ޓ����E�tg��i���aQ(7r���k������@0:��=��P�lC��^�FI�!<7 _��`�Ђ����-8"�#~�_-�j�C=�уҬ�?�|B#:P�-��7#����Jp^J�MCI�Н;�=$��-4f�P�l�RG#�ڹcɶ����f��@�n2p��e�S��9zy�2�p������D�ME j]���x�����ZG��5����ᵗ5q�70(o"��z��d0'^T/�ekt���f����3���ը7F�3�T������	��
�ڙܺ�v��>�����W'��?u6�t�J�ky �X�(;�s�r��3��g��،�y��K�1T+}/2�t�q �v�Q���T+��p4�	�����]{�+Gy1�p���R�ނ�d�ep�\MR��@�d��I�����֧��oI�xl	B��6 �O���;��\B�_uH������bع��_�2β22��ȝ�ۡ��\�F�\W�����7ʀfN�BO�/�i��3��t��Z:��n��j��tC��.��@�P��.0�4$ӛ,��Ȱ���6/�^��k��鉚��x����ʌt�UI�S8,�V���i-��V/L4��A�;�(�gs�#7e�ȅ�ye�8W+�꥜/�_$�[�����oVg�Kh]9�=Z���2�%h����b�}Ώ�o9�ղ8�υ��*O�����_d��$�23�iT�`A��
s�?�X�Ҧ�������$-\��n�2E�ʱ��Cszㄥ��as�pRF���^:�	8���[Q]����o�	���G|�I�K��	'IBK���P�^��0ٟ���jټ:��i�x��1�V�G��Ȍ�Φ¶��jc��ن9��2��o?���D)_�߻��L@��~��^��3ԝ�鬗��B�#�$�c8��.q]n��0�0���,���
�a����wO+�T^�0�-ۥ5+�񰇫H�������c
N;LM����Og�H�ɀ��\G.[���CY$�hP��ϪK���*�Et�G��9��R��5J�h�ى�J�U��I&zVu�p<��K�B�[�@[�������X���;�T ~�����'����WO��2wu5w��e?�2
x���dz)v�}1�8�z�nX�PЧՍ�U��16	�R�J�/`f���Dۗ6b
#O�a��߮Y�
����\a=ݧo�j�?Z&���T�D���|��Y��P�F$ N���'����y��z?U���9�#�Ʉ��hX���9n��,�&�h���]���Z���YM@��h�k��3(���Q�v���7�^�@���>"e�aL�H�{���y��1T�o���/03�Eg��RN�~�]��m*̛�(v+h�چ�-!4I=p ��=�G�,�(�T&��<ߋ�Œ&�Rf8}r��aeh3Gs��������j�1':ͽ�]�5�d���qM�Dd]:����{j(�3�n"�D?5�rT�!��h� ��r����a)��O
ڈ1��o�1D��d5eg�d��_�GK�dU�E(	>���65,Rr�N1�62�;2ol\�k)1w��kI,Y����٠�4l�[jʅ�������h!h�b�y�'��0�����:n��w�,bzK �