XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��_���?�4�4��R�(��O+�x���y6��v�ಲ8��Z/�6�xmT	�2�WZ��D�6*���aڝ�K��.��*�����ߠ�Ä���G$ė�N���c����>���N6GM,Z��O�����%��܏��.{s�I���jȨ�X�)*������W�GG��)?*|Ԭg�԰T#��\;�U�)̏1�1�P�����%���}�k_����$�y�!D�`e��\����ɚ(>�_i��p/�����O�a�gm�Jv��_z��C��ٝ���IO��4�w)�[d) ��^�|{��	��F� �
IQ�-aVo�a[���	�T8�Q����oC��P	j�7�O�Ď��n챚L�L����q�g��/��+ɀ��"�5�`:����tt��͵h���?y�!�������K՘6�g-�î���Ӑ�M$�٣�K���U�b?����+�|l���=7�J�y��6���I����V?����v���A_���OS�����n�Bڮ	0��m�}��:t(W���_�z_z���}	b���}0��Baf��d�,*�~�U�ҋ��O�;,�@��y�Oh�pIm!��I}}��M��,�DX��Ҵ��pbN��E�F�8�R�t�ܽ�|`	W�ZW��qh��?QZ�?����B٦l5�n�`��H��h�g2���0�c2��W�D#Z�_╬ל�rb*35|yK�i�����cd�l'O�0p-��W��$@C���F}�unXlxVHYEB    20bd     a50���
��o���4�b���nʜ�J�X��HK:ۦ>�#h4�$����E`�sr�_���~�yk��Y��~�Vh�@;@�Jz����!�{T�1����N�1�qk�kA�č� +ݨ:����dw!�����!x�?���4ucR�n?'�(K�յ���9�Ǔ��*X��L�2�L4p*���wX6�0�	�(��*�D��74D�(���s��K�L7w�1?x�FUզ'=s{�Tn�	 �$L;�B����+�z��������W.�cL�k2Q�zUUj}+>O�(����>p#�z�:eY�w �A�Jnȷ���e�(�O���{Ic���
0K������Z��s/^�~�~ˏHQ���QBiCM
��'<�O�gqU�poO �b�?(1�۸i�хDj,��Vܸ��q3��_�ත�Fl$�1ȷ]5mh�xW n[d6�(�i������\�B�<��x#�U�>�1$#�����q=�}E�����[��\���|[FW�O��>3��Aa�� �K���;��	pb�%4����5bY��dt#KQ�i�"kț;B��Lƾ�ޥ$�O��x(f��c���$d��^�P	�I�b��W!H���.�����Hs\X96բ^��S����]�E�O)F�+��β����K�#���;f�<�������Ѩ�?��G��<�gqy�i>�{���x�<�_9VęNV��T��z`5j��Ɗ�U�{�s(����p����t�8�X�0rp����)ZZT{��ZPZ�W��C0#���	e.���PP����S륓zr�6p���C��+WkuYЛ���vSs ?�ɿ��Y����Ò��Rf|���+�� �"�K�Q!�����MbǤ[gKPaE����k`j�:~�f#�;���c�΋A�������n�y�l�v9�s�0;i��l4;�u�ɦ4� ��F���Eϝ���@J�t���+��*��(����0��|2�NRt��ȍ�,	�&��d�d�������,=��P��z�ZBb�_���VP��lg�tM��9:z�v*\
M0]/n�j�X���Gⴶ<�����&�H`0�DE��h餲6��r)�@�b��t]Q�N�C����/_GD��Ai��oH��v��g��V4����D�/���B�:���U�e�BL7�K�z9.��>�������ȣն�\���|�9�,%X+Έ�k�E�-)�$�:܁Se�˂�l���#�XO�w�#�$���zoW�c��f�܅��L���k
9[v�������,��Q'�۽f�f��h�R)˄If�x��?�@�3�`(ો
>y�o�k�$����61��$y6�o�Kߢ٬s:�DwkZ�<F�bW�D�s����&����8`��Ny���?�r6+�iJ[v�΁�=���5J���uP�`2�u�lR��ي;�bΠO�tw�������*�̽ӧ|n�h\�� �<�X/y {�j��b��~������)3I�f#�Lȥ3 ���]ޢ���׽Y�N���DH�٫0�����HԴ����>Z!Y�Fگ���8_]�chq_6U_���~������
(��o[{֫V�9�ۭ3�_mRnQ���V͑�͏�U�/K+K�ɘ����bl��;Vb����H�GR��K�r��	z  ô����7?�[_��X�ݘ��B��Y���ʂ��i�z�o����?�`��a�7��B�4�-�ˤ�� �٦����ӓ���{��J�oB���@z���j�T����~����>۾R��>/wp��)�;#���9%������CSX��3?�d�-�~�z�8�s��b>�1[%�A��:� ���Ko���B����?η���o�� d"Z�7-��?D�X��?pń�l�Ujl0qW��Ti���o��1u��#�@|����X�����t��?['��Vu��]��آI�����RM�x�|��l�9����[���Z"�S��պ�Ճ�
+u�c ]q��B��e@�#�5��a�s�d,��Ppqrӹ���eB@���2c�].q��� =�L��$���$�"$N�N30iG�u[��h�b���f��g�L����z�'m�^wD�~	��]�I ~@n��O�mX?��xm�O��q���:����c�l��7���p:�����:�#b����ND�ˌR�]�<�[$�:V|�T���(݁��|�ɣ\�h��y��������c��TT�V�?�e�s|���=�`K�z.�Ř�p�����u��G2&�͵�Hd�U^��ϭ{����qyeK�71O:`���kƀ�Ӻi�����>tz����m��?��20L��"$�)�!������=Ϧ���Y�O��)��.�A\`�"';��M��t��kZ��.�P��ʱ��e�,�[d��:��*��j�S��R2�TL��+��x��!����W�I��t��^�����!��Q;���@���G�s����Y�'	M@e��8�WMr}�;SoAB�z�0�P+SaueR�!�
�٢^^K�n��@㎇+B��H-�_��Ҧ�,�z���10��	�U� �E�b��=�"