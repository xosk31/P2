XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��`��#��ldIq��+����)��J�iB�MC�\Ј��.!Ϫ2��mԹfn(4� ���휞���Ԡ�<Rm^ޫ��d������_'��c/ChW����b��޸�Y�C���]3�[�k+d$�{u�nBYM LA?���(i���h6�J�yO�V+{ւ��:{�:4(G:1_J���Le��;��?��n�ߣ���:�����\�OO#5�/.Na�~22�3�Y�Z��sz���:����\��m�7�Z4׋M�c�*���H��b�� }3`�0sF�o*�o޶C������J]��0�?�DU�'���I�v�&����S�jǫ��;���r��)h
����"/3 �V7�s�c�ybRc��-q�������8�j{ÀX%��JE�1���_.=ۼ��^�8.������E�򌷘�`��6%��u�%Č��������XI��j� B�V��� Z���Ή-�}M����9}�O��̩�9� ���"�1Y�H�u7��&!"+$6P(�B��	M�� `��s�O>˨[�������wLF�b�o�#[u����c�-�t)��lp7�ʺ����$�x�y��j����7�p��E!�3:�`����&���q�Ϊ���"�ged���O�[m�`3��<C#�#.[�!k�i�����2�б�����YLkaI1�c\:im�_`��s�Q�{s#c_]l�s�u�����~�a
�}�
"�l籱����rM�-,����<2h�Ֆ�Ǉ3I[��{�]-Nʻ��XlxVHYEB    77d6    16f0[����F���W	����L�^�s^G#�4�'��[/8��aC�M����րefTpW����:BR�5��H�ꏀ�<�r�@֞�t�q��g%
�=Ў�2u?O)�]yW㳛�ST�k����
����B�$
6_��"3���-6&�fV6%�7�p#��64��wӅ_0:VA:mb�'�^����L�|�':�Ҟ�עe�/�2��s#�	����%�2c����.*��%J~��48}׉Dv�)���Qp���|99��!�1nJj}�xʍW7�[�ʗk�Α��cS�Y��	�g@��v�p@��d��'-9���Q!��ӃF$�:�����oZeK�5�+��:�(��C{�ԁo�$��g�p�/{]���.����B!��s>o��o�܍�I�Y���l+˕�;���k���~ {��� ��T� �y�>
[�g"v�c��j�����~�l|.v�jA,�ʽ],�ö���VL�wpj�5tD�vr��s�wؕ�g���m�����8�	t��hr�}��&kpؐOm��@#�5����-�2��1��rI������Y��77��!t�_VX,�%ǝ��}!�3؍�M9B�_l�/¢=}���1Di���C<&���Pg?V�
@��=.��H1�a)�E��CyU.���G�1ܙ�6�a��#�j,���ץ�#%��9e!�!�~�&�|�r΍Ϸ�9T�Ό{]�j�4
m���KW6��o��Y�����K�i�.ܖ�v��yc#[l�L�g��P��yXY��SI3� �i�:�Y��,$���L7O���]@Àݏ�RaT�znj��`T� ���D/�Q�>+䶭�B%�Sb�W�}p�����Flv��ӿA<y��cV��[�-Ara R$Z6)�Ȼ�d7�Ji���32\����'S��
���2'���_�x��x��i��7,3z�b�ϫ���zZ�qE����k���W�cK+��(o`w���jfj�9�Ȇ��g�
n���B�[���T����>�U��Y����Xb�u;��3幖��re ~�	O1&q�չ����KQQx/�׃�؆��Oȶ��#��"�ߕ�*��YZ�[�R)������[����<}n�&F�������<��Ev�g(oqb���2���D?�ᱳ=�+^}���PeT&p7 J+�o�l�Q_�=���!D�}�q5��O�p��LK�͌4r������[Wo\TL(A҇<��i7�d���e�%�R&��,���������>�q;��L��U�R	�P)|��R�+ƞ5��!(��ؿ��OV�W�/�ki��1�
LJ U���3�.[�d�O��(�"=R����\�F�ykϳ���N��)>Lsy��3O �ލ�$JV�߲~|�ީ���ud ������s�3�K,>-�|Y����� �E��	.��_��h}1��:�U���#��rp����j����n��nݫ�b��I2�����tx�ˋ�Y��H��q&�8RW|�G�̗T[OeB�4�UcKB��� }����#67C����hS�p���99E\V��2�W`@� ��m�!�->��X��U���J��O	
$���e\�V���|3���ok)��AԢ���>e��`P�z�Æ`e$A����(F1(��!�I���ě
"(;�mVl��4=%9�c?lG� �Q�,/>F�5ߊw�:�%����
����[N��J*/��Ȩ� ������S�YdV���h|;�h{ ���!�Yh/�h�B�K��"p�
�W��%�/Bծ���}2��sس'a�:�\��ڢ�A��������pZ�^!9xG�M�_{�O�uN�~��s�+/��1v�q�b�r�Fd�5"Fi���\a'���p���`��$���8N,P�x]"ʼ������
y��پP��L�����>��7Y�[{ I<�wm��gPjg��.F`��* ��+�x���LG�� 7��	od	���H���%ߊZ^���,����$��"<S���d�R��Qg2���D,
K�y�s����M�m�O���������_�m�V��$�0曺��N��f�/8L)��q��,�)uAW�p�f18��O~e���҉aE���8 ��2�,؝E�_��1��j<)���t6�$c��:�L%�ѿ����������E͔��ۜ�c{��F2l}L��X�e@h��"$^��D�J7���4'"��� �l��2@ (��QE�i�"��5>8UUc[�._�_�i�(o3�߂�������h�mģ��Iec*_3��֑�>�֕��!���R�f�&�:h�cP�Қe"�hb7+�k���rMHk�Z�s�^`tW�ID�4���^��Y2a��]����"�_�d�ޝZ��Hሎ'\$;zLyA��]��0�f!�۪jɐLi~r�R%2�>(O$=�{]>��&D����cV��R���#qҤ�)����~�K���G�g��o�\G�
��� Y���,� ܡ^�����l�.f��q�Y۝�p� I��/�������y�r���W8��Hi��yR�G2<wG6�Z��3O��iqjkm�d����,��Φ(�9hy��d��ٶ~�$��Fy2��|�VsW����W�����궄��~�v4��j��L5�p��%����	G�т��k��ъq��ɸ�C�
ܴQ��<���_�z���Kw����X���|���g�#��f[[��;wBKٶ�g�6({����,���ц� Gq�h����+��(�0��#�V��<���W�s)�{�,�+�����'��h#�m�'"�8��ԃ��<�_�V��;^[?�BS ŋ���~
���ύ�^�Fh|�����.-z��~���î�駱�T�!%��~ 沅!���Tkr�ǲ�r�5� �Ϯ�0�;��7p�����$jY��Beg"���lY���,ɼ?�d'7o��v���ȟ�_?�!)_�MI�9���B��]��Bf5�+�!I�k&^q��q��s͹���Wm�GҴɛي�ZG�>��u �xN�*��)cq4��A͚͟�{�����A�� �'��Z��E�3��+߀z�d������wNŶ�2^�ێt@f��/����$��1-N�����]�Y&��G���~�RSg�u�-"��e	x�t�$z%�Xq
"��z����1IK���a7]�T!l3���f�$�:��K��wk��H�S�S7z��"���_1�O��L��������T+ԡS�/�T��~�3���|�ާNڏ��+�E���v��`<cT�(H�hL�(j��#$Zr�4��K��?O��vʢ��١��3��SL����PR��1�4۞�c�l�]�������)p�^�h�N�B 0;�?�,�"O�j%o�88��9G��\�8�֎2.��q���
\{=,O�kf\���O%=):1���SoY(J��i~󴤩����k����θ�����#��V
�+6�J�=�㩜���I���3�=/�Ŭq^E��#�q|��M�˃$SzzG����n���\�����
[��(�(ʌ2\���ݝ1R�6�'�K	Ҽ]Q�k����_���	�ޥ>�YXu�3�n罋0x(�f�D�z?�k6=Y��]�`P_� )0~k��� ��N��$L���\z��(�_�d՞�y���6���'b�m��=e-G��Z��E�nǃ�25��t��M�a�� &G�-$�6�K~8��5�iMN����c��]%��,}z(�ܲ0�z&&	�2��M�<;=�	�����܈O�Q����;X�N�xN�|ݓ-5||П�7�?R�a�냒�j&T�"��f��Q�OE�y0B�$ޓ�(�{z���՞?:+'�r��{���֍*�>���i=�B�ǥ�z�t�D7���v� � �FY|�HM�9�Ȍ�Ͽ���
���ٔ{-�nV�s�Pl��Ɋ�M��R�ŧD��5p(ص�ӌ8��6�
(��e���U�>kJ_A�Mc�_�� 6uXr՗�II����(�0�uk8�_I���T��W*@[��?B��b|��l��]�hIay;S�F�Qjv���C�Riu����r(��&��`�߰Tn�����0ṷ��>�����q�* r�/*aR��"
�.ҷ���0��yI*c	�b� �d�8��՜��b�ˣ����~S75s*ژ��|�D�����s9�/����z��J0���Zl�Mv0*�r�].#p�∙�+]��w�%��Xd}G����)�����M�+X+W��>�E�a��>�`�[h���%F3����JS?@@g�F�x�T��3��㽛���@3]��������M}�ln�s���!�n0�g�{!��5y.О^�v!�m���t�b���r��O�	��@%<������1E��0jZ�Dl�ھ��O�d�է�y<T�٥@0��������[2g|M&��	� �ł�j���W�Y��0\M"�f�Q�������)��ɶD����)�=�?H��qҩ(Ⱦ�N����W��B�m��v�).}�K���32<PݘP�߹^�SX���B��������aX��d�k����h/,�wU��I����''&�z!�tx���^���*�BN�%Wu�m��/(ؚ }ߊ��4��K��7@k?�#��'�n)��#*21�̕�q�ड़~��m6
Mڴ����ZVbF�O� ��ɍ�읫I�X�m6:2X��]�7�=�F�(��N���Đ�/� �	FVX41l��LK�j��q�T�����l8��՛�r��_��Ztx������OY�.���K�NǦ��S�e�e�H���S���>�����D�c�|�f��s͟*·;t/��B�R�n��x�S~�[�����C��*��l����p�6�� �z�SЦ��5�gIs7y�'2����MhbÎT�E�LQ+�_��&!��~ĭ�2�����3���F�5�2"��w�J ��N�Lؙ�� Y��>ظ���vq��#�P�� ���?'�'�	<b���:����/[��Ͼ��=�	Ӱ;�Wc �Z��%�y���k)^���m�#2�e��P8��5��;�g-� MS�B	��9^����,�q"{x
�Dk��� G�}�����4v��=��*�ȓ[<��Gp�Q������&�ȍ^W�;��,��}��Ok_���P�l�q/ �gָ��ׁx�Ӯ���}z�p&��=���E�t����- �p��ZuWp��H�i��=���R��'�&���<, )%�`���i�x�Q�֣�E���!���s��Ul9��1٪��&7 Ks�{j�Gc�����"��߳���Q��6ߘ�����s��J]��i�L���
�(����!�109�{�z3��]��q#�@�/wi��D�A�_� ;��uzɐ3��Ud��Z����V�@13.�*�T���XM�d(��Ē��q�N��X�Ei]��g<��wҍA�ͳ���V�l
\�.���d��e�e@$���J!b���-��F�`�2���\�$��|�a���}$L����5c���_>9�`��9\��?��ɝEb�I1	�����D����*�!&:� �e8΃<q�<WY��p�	�J��?K�D��O�"wRY*@��>����k>�T(�����+����|�j��gc�Fr�S��dt��q�a�~^�R�� ~����氙��'J+�DI_F����:�Q�FC���Jn����%5��+?