XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��5V%x��`�a��K�TJΩ}J��p�J��!({�%��$�wF�*-^^􌦳�����>N��S����l	�]�P\3*r	ug��1�������?��F,c
%�㠜i����Ҡ���^���(���+�6#]e�=!���,o�ֆ���P�1�3�.��/wy�o�ٚ��\��88��|�Յ��K��vbQ;��m��ޞF�۽��Ȗ��;�,�i:��B$����)����,/�Pa�=�tH���K	Qn���r'�*����*�������,�cq�Gݗ�1�U�:�r}��7�%)q��d��YM7�Ol��Kk��E��Z���F�_�O���Kص����	5�d	;��AZ���a�����9��.�)�<X�q�7i��֫">4V�J=���C�����LH����+k�-o��eB?��>ơ�B�՜�^�F�KEO�� ╄��in�E������^��#��]���
!Jn:Sv��gN16�A��`B�h#�û7K���>�����o���9���X���1`���M\�]#�`7/�P��әj��S;\6	s��[���D^:��%���0yu�K�d��n�ijc����x[u]�V3��'(}�~:5���n�w�m'��?��A0��M�8�]�:~&�O{���QDh�d�Z5F!��}������5�.{�U2�&�f8c�!w�f���Dʸ^}���H���կZ���\35��v��Ie�\�?<���B(�t61³�XlxVHYEB    5073    1100O֧;��[�L�sM����,?I�C��}���65\�А�(�(m��t���Dd�����p��@�`�+B::|��͹�T�,��D�3�V��b�_��:Q�gv�+�z���,����Ԡ��{GY	����/Ӓ��t�!�E] �:�Ɨs��,��ՃC�����_�u�78A��,Q�q����St_^�q��N��qF#t����|�z�fr�	ܞ�7*L�=]>�2Y�F3m[�J����=�Ŀ��DV%�r��#��b�!���Mv�Ax���k߬VV>����K�,��q�0�Q�$m����2�J�G�Ne�4����x�1����}�<���^ї�=������
��Xp)[�)�Ǻ��[�0�8~���$!V��Ĺ� v��]�<�Lw��#�'	s"��{�):O����$s�:=N1��z�5/����18X����a>�R��x��m#�4�����7N� ���ǣCp��ӕ4��e"}�]�ƙ`����P�>j�l
r�o��GEw����t�c�T8��z�m�r�Ua��Wj~��,��e�*\��X����e���CP"`BK��V�h�`���AtJ���<굿�i�~�$5���?�_z��u��	|5ܫb�,\%=¼�i�k�Ms��#�X�B�O��'a�Yf�7\�g��|����%9�B0�r:5��j�J%��xq�G�������%�j&E�B��@W(��0ߤt�P� �x�-�Iҿ,���A�����*ߧ�~��|��l�u?-ɟ7{�!��d�mx��.���+�rx��PKRG@�ߢ*�_b���+M�6���3�����!���Y�����J	o� R��as%�n�SYf���s�]&�nT1P�6)���apDCp��oP�6K�'��Au蔦n�@�/3iM?�w1����I������).+q+.A�o
�w :Q�5�K<��L��'��є��X��� Y�W�����	]����]"#�1���jt6����,�R68�?k�)�@ڽ�< �~K��3#���w��k��D\�Z><!{I�	$;17-�4Q�j�lz�*���<��#��
�0����R����\�P�N]�4cڄ�h�B-��c��xNv���9���>}`�kt��"~3̚�5G'��tHV�� ���e�<�����x��P����t��<k�g*���ZȐ�%pAO��6��u�aH{�:d�,��1�~1��+�X���=�Y���)��:c�E��KR���s�Vkp��|<	�Rܲ}�"����Pq�����.�-�[7����YY�:/ز��N�0U�ΆK���,�������� ���u�aA0�X�F�ge�I�1�O����o�>��˶�i#׳X�	��̸5�f��M��{�-cK��l�o�A2�-����o
C���	���0��JV��ず��<p^��-\W�G��%S�уc�ϳk��1�T��_�@�*P���)�W�>3$�;m���� 9�<�����"m�n�G.A�)�[t�H*zAN�;e��8*U�)�/_+P����#�=S�)#�ɗ�� 4�<R@.��*gw�76l� �R��b��4W�bG�R�W=�}ă���5~~�-i��yN��5C�T�f�7e�e�Ӂ9�l5,�x�S��s�T&�߯%�ɤ�n��8��K:���y%���!	k"�[���ؒ���OJ����]/	nSk%��d˦��\��
�3�S�#�.�4ڏ���U9���Eh��΅܌��A���[�jהp)Cy�rj4���<�����P��WǮ��G�n�ڿ-{��K��)Â�R�G�( ��H�Uc��Ì�
�Z��S�=&��'��8�\���������+��]6X/=b`��>��a�>����Y��WچG�s���X&uBGPS�R���7�9���=�\�xS6x�<�(c�h�;�c=?�)��Y��x#�[$�u�����*���la]���/�9N�`qXq�g� ��Y�3٨[K��Ca��������W2��f�f\�4�k�޳������&�+,�Yb�؊���϶J��4�<w�&NJ����H��/��W�����x��C^3�$~e�������2WL����j(h��+�
���z��$����N��&�D䠅�=���;"1�o�F R0��I0�/��.E@[#n%��\t)O,�e���T�Zd��gM��hu�sn���{^�rC�o
�� ����:0e۔[p�V����֖{�����g�^�[V.y¹��!\�T�p**�����Pݼ���χ�s�W
㢭l�KO�_Yg�:#,6�?U��\����Yk�)ZFf�0 �NB���@;�D�#��n�㨚���}i�����/<�i%�o8���z��B�^�8Ti����M��k�{`��,�
�p�D�E`2,]咛K�B_�:	)��@sŵ��U
e�l�������b@� ^���r�����I�]!�i)�s��#FC��ҵ�ؗ��$<]Xп�I � F�&� �Kk1k�R���A���]VѶ�������'F��ot���<�Ն���$�_�}������I��F~�+9��c_7sl�Vg�6�@D̯4{D�,�Z.���Dz��N��K�F���������0�ٿh�f�<�]�~��?k7�08�o��-��*��McQ�q������P1��=0��q�BM�:&�w���f�լ����^n[��	*��C͒ud6~� �Q]�.��mE����O����������mpF�~8u�I�ڟn!Yy+�ֵ��Z�!\>W΄���pi�%^�$4�C�9B e�&3���J$�o�;g!8iMM�s�=�A�i��E�����Tb)	��|O����P3�,�'v����Ą��@���>o�~C�ͤ�6�u��Ǡ�q���,sB�gq�]3fI����])+2
:4�#�IH��OiDx�iHK6o��{��Mt�����/
�s�ʟ��$c�_70&�RG*f�J�1��\X�X��]U
�0cP�2� ���@��xH�(�Q��~�ܑ�9y+yl�JG�S<����Q!����<�b'�x��m#�L�����9�����7�.'�n����YH�Siu׿��?�F��H�3�G�o	G�T����/ �^��8;�u>W/���CtG A��|��N�)�"ܷ�i���#�)�6�\{���Yc�w�g��o�f�&�w��������y�@T4�L�xO��d��Eb��/ƂW��u���_���u���İ`��Қ]�ntч�v�0��-������Gg��4����w�r���L��uY�[��T_DGٳD�/8@�h슼e;t�����`TBne����0D�Xqv��A�+�n5q�����=��W��qg�f������T3E $���v0��K�<>�����$�D�h*�=x)!����7�uˬ���^�14���l<�c����*���*{'�YD�*ę�����ڙ�~�'r��_�J��Į��ǿ�Jڙ4um_2!�4�ž&����Vi4'BK3��;[�LI�m�Y]�X���=&�:�=��KN����|�lc�Q����&,�� �r�rh�t<�������.�x:#	�q��>�e�y��F@�ew�U���� f1�ND���e�rG�0��KB{2c���	=��0ûC`�X��y�"Ej��A`��[��5\s8�u�#^d�;��^�S,>��#`��M㒳ː�h�����x�|.J��#���-���4�ٟζ�=8����@�+��^�];Ј���:�T�[���CWeD�c ��#f.�\�)���b�cD�3w�vpՄ9&IwY�_�Cm��`.���M��/���WF�V���[Q�	�
	�-���������0�L����5����� X
XF"�LA����/�$�1n:Gӟv���w�%ľ5Hp�s�)�$7�r��6b��K��GL���_X�;:�K�H*a�����rݠxݨ��[n��q_räxR���%�
;bm����׎�{����%�N.��rA���M=>�=��N)�������r��W�'�z�̑�׍̂����SH<��N��#��܏�+�0�_`*v�@�KT��G(�:RP��z0��H�٩�Ih�D���-�����F��Dz�-��ܝRQU�%6��+e+)8�����q�Wؔ�gG�R2nYF��?'V�N؍zm