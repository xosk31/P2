XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���+�����N%��p��OkE5�6��Y�)�VP4X�ʈ��ݤ�1��~_JLۜΆ��.��$,J8���t��@AFa6n�%^��D8�2�v��~D��_!z��ҥ;�A{����Gcܣ���8�%H&KI}����wAN��\6;W�g��cUR> D���	��8�l($pI�}ƪ�^S!�Ϋ>�9ZcBp���V��r&���D�w�jʖ������Z�5'81�x�5�V;D:;�;3�W��@�	�FB�-��7��[e6�I���1/V$�av�I&[�qeQ<O����|潦���*0�1�@q*�=�,���n�H�#�'���z��A�'�s�'ĥ�m8��z�cr��1'�:�<�q~���]Q����P��4�O�px��7ϕA	b���h��	��I7�R��~<F��C���%[5��4_�+���c��f����$�8�)2Lr%�O�%������Y��6
[j�zʋk�����H�eS+�|c�(�"C��jG���k�����7�d1j��:!�x�1U��U�N��3�Z�����W�Y�a-1��-�7k�"����-�/H�G��s1��A9t-3�ȓ*FC������� ����i��P�������~�I���$�C𼁩e��/�Y�V�f��st��Ǫ?����&�ߗ��J�b�Yj��a�nIۂ��,,���A
F�� ��o��s����r��s��)��o��� A�<�l�SV7�Q�b	��_q��V�XlxVHYEB    fa00    2480x����(3��MdV���a7	v�o(ք����D���>R{�qN6~ӌ���'���J{$-!�#�N�l"`\ﵳh�_9�p�PB����O٪ �S�}�* wb�]���vi䵃R�q�y�q�������W�k�#�H��cޟ�o�@���93v4��ޕ�nN���^�Z�b��B�O�9	8�ELޑ�Y��r�I�S�`�4۰�HtV�Ү�ZE�� ~xؗw�MKe:^l���F`�c���;�UN4��
u�ޣ�������
}�B��:}�=1���^����-��+��}Td~�]m=�藱%�{(hc�쵝75�/�Dِ���R��征�ı0���Č�R��b�{*؆�[W1�����z�.?I�G��q�
5��lz�5�%Fq������JF{�i���,�<�R��1>.?a��-��x���ø�\���+N?{�T{��y�n$�ۦ��
Pk�^;C�*�L�f��狰�F4 ~��8]��zX0���fF5���45W� E��g*���m �U�g6!��'��K���I���@	�+�LY�"�W���Zg��q�b�����Ż�%�F,x�&�E�ex��V#��d�DO~�B�M�d�<��A�n�%����|�U��ҫh-'��Yyz�n�G�&�� �f���Y�&�� �S�Q[~H�	��<0gD�ZտhΞ(�f낤b�S����ϔ|*n}L��*"C���8�-�秩��J�G�*�ߩnfw�^����ݎ>���:�=�r`p�yYl��Q���Zg4xD
[$�l��N��PMb�
B�
0�#�5_v�ֿuA��D�I�o��Q�9�l�v�?J��T!��j^4�	w$���anG�d��`��C���b��ߚ�H�{�N�Bjnv%]�=)����q0�ª�Lh-2�����G��S����Jh���j�'�l���8dԚKԁ����ԣ�iEǵ..�:+��JHn�B/G2����+����]�0Nv���c��c9��[O���"�'�6ZW��C#\�	?�k��j���%A��t�*�_<;-q�7����,�E�
' }�>��**���[��G�E�}\󨌌��߆JsX�?�Q����F��Ҭ�QL�܈J�)<��S�e�����]W&*/����*~�5�jA�_L�G-�����ˆ�ǭ�d̠�O½�蠱��W��,�:0^:6�1]�z{ocN�FQ�b�EE5J/,�ڟ��(R�W�n>�S3a}�l�`�뙛
��t��S
'ފ�\���}�R�G�_��(�TT����=�8��G�c��w�j���I�Y�ɓ�bCzq�V鱆^���P#�Pv�f.��5��tl�R��HP(��\0��|�����uD�Ǵ	1�]W��n<z��yc1V0=��,�%��&�ۨ.@=�78�:�_����l�~ �FL�6>-��~D����7`Z�D�&�O.��.s�>��Am�E��F8"�
�O��r��g�PJ2�WO��32�k}=O�q�����WK��8�$)zb!߹Ác~��ƖgǪ=μ���@3����ׅ}�r&s���a�*mk�Q̈́I��=7����0o�~E���K��1��g��n���)g@3��J�����ۀqu6x�W�q]��H��ʀ�����:�o��.�<b
	���K/u�[k�@9��I�cva-M��ED��zi�ȋk\y5Tn{���Cy4���8ۛ�?�c�K)�7!��\��>�S�&N|���9��ߜ������=�Z�%�N^��$t�Ӿ��;�h)t���@	*�Ix���T�8E�tMM�z���t#�ɋ��gb%��fӳ����6���ҭ0d���U��CR�������)i�*�S �p���J��ik�>Ҋ����f��� "M��2�Yi�<�f0��w�g��a�c]�S5��<R���4��u�&��K�|�*x<�������	���(:~�Fy��-�3#�4�ދA�}_e%3w�rQlL&&'C�tC����-�P`�?|��u���&��2�IU��&7cw���a5��?�N���_�IQ�����!��j $�C���#�Iܙ����@� ��CѪ��l�����%�h� `p��X�t����h�1�ʘ?�@>O���).������5ON���_&ȏ�8Z��eRu�$J�R�4b�؛��� fڪ{�{�{^�fT�R�Ee�a P?$��zk�.��/�5����Te���ɮ0���yr}���9e-|Z3T��"<�m�lS�o�s\�ZD/���/F���~��$���.��C񐐀�$��}���^�v۫�͙@���.�p����S48?�N#�X@_��S{�#���J�P'�7�=�,���F��`&�����H���m�F�i4]Ϲx���&�
F�<�^����2!�,`��h����KC��{qwiG�F��<���~  �P���2VM t^״C�i�o�/�,�U�y�d�M�`	}�K�(�w��$��:��o�X�P=�V�Ž�ꏕp��j�p�@�T�:�d�}C��Ԥ���e!{�P�M� 7��粠�-�6^t��������7"��c�/"WU��4���#�c�V��l���'#^��=�,��;�h�~Ew�&Y�y�TK�2���)2�MK�vEGzf4q��e�%��G>9�F4�"}X>��Uy�J�PY��}UQ֧1'�_|'k�T�(6���ͤ���)�!�"�5W��I�ٜ��s!���=_> ��
��F�j�	>��E��i
�X��4+�}
���ɐd�Kh�W�B��H�Ӫ�6����,���1A��K7��9�5����@�(�p�zR���d�O��i4���P�x��K>HM�ь�*
	��,�TA+������d*XC/Y�R�%�k2���g8�Q�(�+N��l{��\��V�D�=i���WJ�&����I�;⪢?&g�1~�M����p՟��+��ۦ�2�%%~K��}�vB�TGZT�˳�L��ފ¢���"��9�bM&������[�#����>��"<2PL=2�gU�wż��&Ak����y�v#w�)�K �n�:���Xz3_��q�-��+���	�/���1e���ʪF�F
���߈1��X��Mn�ɪ]v,�}WK3���C:�G}�+$^��-E�*�>B�~?���
Z��a�n�N�����k8�t/�OYo�e�ئ�����=����Wo��f�<�(�a��$�'�3����8�����y?�I�Ϊh+�&"An�����}ΐ�\Fn��5�!\��J�e`a693扢�>B��_����k��~F�VBC5�ʩ10iq�����@F[��.�E�pz�I�S�d�Zc���"?�N�=y�8��q�}�B��t
a*��a��+�*��N:�\�����
�HA�d���k�7�)Vtoq���%A+��S2c�S4AӐ�ݿ���L��]%{��EXM�7�_`�,�7�9���Ʀ�>�����lDa��.j����y�
����Dag�)�m?�/ě��dB5e�o���1F��W<n���a���S�bQ؇�j�ug��W���HF����+6,��dH�D���CIsߟ�)�z�4^��,�)�a¨T�ɘJ���6B*K�T��Jk{����n((����V5}��2���ϛ���sU��M��{�MC���+���#�No��p�Ы��ٯO&� W-;��@b��ہCʒC�Vv�t[L�^�d���Q��w��M5�֟742���`�q�d�d����ڨ*`�	=��r͙�.�҉�2�nH�wIA�z������W�/��mO�.�Oܚ~�⋲/ro<4<�]����2]>�OvWr��jEGx��4� �X��4��6��fYhhq������@d	�4��j�3�W�^�7	<�bF��s�V� �Hõ�>��p�O���f�/�@�3�����M����/4	g.�����ffh?|b����R�����tJ��,�ֵ_�S��v8z�*�h���!�����`���7-'�/^��>k�0�}F���mM�'��a�r4R �����ƍ��x�:A���S:F���/x|VO�r7�CI��ؘɿ��G'ӽ��y���M�4)��E}�x��4��Ǜ:*��C�U��He�]����������b:aYN�{��EUCY5`A�y~	T�/kҺk��5%C�w_�u�X�W����d�����;��0��#���O����1��;a���1�-�Qo.����n�:mZ����X4��vR��j��p1�`=3<�ؒ���~�j�	��xI%Mٝ�����vo�̆��se8 w��9wDY3v�	���l(o9��O¾^�J/#�� s�N��B)r���c��6���Dj0Zk��-��b����:�GWe�O�T�<cTâ�$#�r�*NU ����	�|JO�l�:x���B�C�Sޢ��[I��5A�6�(����~*��V7���t.�<a׾0O%�}�P0Y�=��ze:�S$)�q�E������
�C��2��R�Ӷtv�,A��I(e#o]{�АΘ �v��J]g�pGa�%#����)/�H=�k�Bf�o���� �"�*���.qBzg��CYW�0�N��-��7��y��i{�B���/-��&c��k5�'���^s���L��WU��K;ˎR��P�=&��:_`�x����;������߼֬ݾZv��s�7+��P[��&���P��E�����3��N��J����z�8U����AR��Fn|� ��/M�Qb]q���BQ�G��(&�3�M�h����Z�V�/��sy,�Q���BL��!�I;z-%�9��`[����8W���'h�Bk��:�	��ݧc��������s� sZ_�%���C'J�S-�wVO��tiԂH�,�
�L�
ޔ��f\�q��X��r{�9����Ú�I�����}B�ˉ&���+�8M�8�C,�pN�N����Uܝvw�����G���D�`�ɐ<��/�U�3���؎�W2`Q���
�/��ʌ����Igj�Y}=+&�j�a�!N{	%�4��01�eDC�&e�r#�Yұ��vj�#�'gcY`�[���10*��c4�%��#tsz��,ߧ���m��tv�a�5M5�8�}���w��E�����F�[��n�Gi�`~1|Xwd�L<�p��dnN�v��ϧ\k:��x�t��9��*�]j�D=�����)��H�J�k��v���aƗQ^���.��+�"���2{k�%N��Z_��9b[�-\���2H�]�v��/������4���2{��R�@�L�o�==f��,����z��	��&�p$b{� [����	��XE��b-��Ə�ɏ]��G;�L:鲩�d��Ώ:Z0�����|�}Ⳙi�:�h�Z�n���t���|�j=D�R�뺎�Do����̋rÓ�߁FC
�!c�X?S�$~�De����0��8.��*6�O��S�9�.i�B���$}�ҕ���P�%4&��sq������8Fo� Q����[S�I���p"@��N'�
C�hR�#D��B'3�4֠!��_�T_/�~��,�0j��3Y1mpCl<j��7�t�O�=�p\B,pO:�3*��<>�$]�\��f*��˕p��X-�љ�4�8��>W�<])ł�S�����ђ�m�N9A�z��B�6X;J*Ñ�T����;[���i�|�@��:U���B���!�DB��, G|�ש��ք��(����]���M�m7L��� �cG;�2������v�p9mv~�U]@��0�S$QN�ܪ7�E�H����{� EI�h3��e�Jܬ損Qo����\�$0 �*�<�85Q�M~r��#���=*x�KJGXI���=���Pp�܁�j�KxBӔW+&�M0ٙƎ�lc�ycD��/"~��>2RV�ZHq/{yqn�0x���E������Q�Я!�Q6���j�QY6�J�.��Aw-R�ƭ�6깵������쯔6T�$E�5v�|���N��\̣K���΢L^�y&�.�����N.�I�ú(:��R/(�@�2�?(�f�Ҳ}�228q�w�Nw��/L�sx����xx6=�=__vݞ��͋���(�/d1��0w��.W���4C�g
��gQ��@�!� @; ��*ȕ9Ӌu�AWq�T�I��F���J6�� �~hG�m��_w}����;R�����֧����@�������c"�Ή�ȿ���v�ߵ��s�,��qt�y[&e�LM4���J���p�&Yy�<���\�8ݗA�R�J�����Qs#���$�Tp{	�O�@�K���A��50�I,z�¶�9*<�,m/
�7
Y.է�J�a��V�H|9
�#0�~�2�7�~^�$�,T��k�����e�B!r��x�A�jq���fZ��EVC���#�j?�N0$A��y��1��o��X5/��"�>a"]�=V��l3�4l� ���4n,�����ŽM�B;�ƣ[���\��]�u	���'(P{ Tn!���DR���N���7ƪ�R��ރ��S^�� n�Rwm�+~e6U#�8X��ݽ��F�G���n�6.�N���F�~GD�E�]v!��*��X��[.�������d��R��W ��Cծelf5�y;Π ���FB5��>-!nVD�_��L{�= �J�O����A$⦪>���A^#�'7Z�`��Vq��,>?A����2����1��h����ubWc��h)�W�G^��\ 3��  OX�c��Z��M�A��#ͼv�Z7>p��B������4#�!X�����\��p��Yl|����2	�� ]�k����T`$�f-9'���1t	�0,G���`|\��bb��[����ƀ��
�w;J�����|Yd�l׀%�;n�����=�� >0���R�w����_�(�ѕT�<m�����>� ������UQ1Gj�ʉ%�_�Q���yB��6�q�a��o+=��̉p��X�M7q(7oxB,��yuC�T�|�ïM}�Xs �zm�0�� ����Ꮵ!�� r��a����I��Ϝ�g_�5�a�[���b���5�g/�Q+�lr�E���al�:�d�`�X�q<��@�X�h#�k�E^Sk~�Nc2�]L�ރH�8�����,�SٙZ���d�����C�{���w�G�<$�Ï/CWI��6��:X��%�頶c��5�vim�#ʖ�NV���O�+N3X
��x;�Ą��q��g�{����Պ�uy�-k�L��iT�Q0R�"�dP?�`�|Q���~I|��h��A�H�٠�w��%֠)��9��3��H�Q��o���jE�7��w�u�xd˸P@�rlO1�O���6�%F�B�{� �KP���$)�8��&�['�"��C�3$�u�ۚ���g�wu��g���k���s�!S�������*�h\�rk���Z�WS��=M��1;�>[�%3/�XrTۤY��ɫcJm�s������lJ2R�(�k˾�ۀǾХ��s�q���l��1�Qo���J�����k᳹�Wf�5�^�5�z$j��%�ڰ�U����ߙ/.�Z9���M��n���=`���c��qc���+�N�b�w3�#��s2�p`Db�T� 	C@\��r�6$#�&���[���hFx�AS��.�#2_
�\}�����������y41���VI��6Ϧ߉�i1�iEl �9����N��q��5=���K
�������##>�b��|"��_�2p�u;�I�;V5N��?�Ѓ��)-<���!�"�wǨ
^�	:�_h���or{�u1e��S���#���]�NȘȕ�0���ݓ�b��ʵ���
�ty�N��c�[�	:{��]��@ۻ���� ׻<�p�!07�>,��hzeI+!�hxgI��-*�����~z����ԋ[��V~�ћ\���!~�E���^pDq��frrK�p�zƱ�U��Ax�]�=�{��� ��s.c����qr{PE5�z��"�c���,��i�6 S�D� e�tq=�X�b)ϣ��Z� ��5�oP�m+	��wEr�B��-�c�l�b&�&Y%ߐ��S���,
����h��W��
� d��M]SܲV��C�|cJ�t��2���-'<�U[���@��"�3^>P�?���3�_��e֕�ɰ[s���s���b��SJ1j������I��L��e^��jH��$NEփ���+�-�Q�HMt[g.�YX�b+t~{�y,�å� �Ȃ��^쮃��tN9�ˉ�$+ֺy1��.GFr{�?d������W�^���gh�&���T��;�3��.��aQR�ѕ��W�jF]ǰ�}�q�ZD�D��+��X]պ]����ߪ_�����3|�lw�XjF�Z0��X�z��� �r�"�Mk�Jڠ��^������ǐ�|ǯnv�z��@$�E�%�_֮>�9����E��L�~�O���4���z�, G���u��ZqSLY_�x�ѡ2,��Z�yGs���P[�_J�o\�&��wE��;<?�O�����pFo�ٴ�+;^A�����#?㑭B�6����}j�g&��cM=��?�u�r(���*�X���5 �a?��מ<���������(�v���
�v���j���1.��y^^{u�S\|��|�V����F����t�xΆJ������n>{��[Ւ�QJM�K�|�W i�	�ڗ�JP����e�g;V����=���n�jh�(3�+��}�j��ߩӠ��6��hH�;Ml�OL��0"�dbA*��Y[�S����Yu�O����#�Sχt���nH�z$��e�����%dH5c�4��p �BQ�\��ޔD,�O4��E�_���I�����ꚸ��<�$;%��K��\G��u�o_�=�e%x���\��[,����KK0�U�=����A� �V7D�9D�[��@���<���38�y#�	+�Q�1}�H�ہ��4Aq&��/dR�W��O�;�!j�{D53��^M��Jn�Oy�U�N��)���Ж�	��~	��Y����@��KO��,��A	g�s���एAb��UJV�.�Kʟ���<�B�j�=5��p�!�{z���f;����H2��9��1;!�xI��BeP�&�HXlxVHYEB    964e    1150&���ե��C�`8�IZ�J��KY}��v��o�|cD��􃌯OsoVü��q�^`N����EM-&i;���3i�=��d
��<��|��Mr�b�h�؄,�U]52��P[E���D> ��Z�	"vP��6X��5�֜��@���v;��
�׏�2K���'��kU#&&�G���i���Gs���_7���zb@@Β�F�V1#�����# ���i?t�5��}� uI������	��������z�fAT�j��H�l/���C�y~l���|�ˆcI����+wĲUb�D9kP��t;�PA��ꀋ$J4���Uu���WX�s�� ko^s�|a�[Z��ߗJ�A@Sa��/{^͂�=�Oj���> z��b$�J�-��損���&h�W/��v"ϥ���T!�>�����x�:G�,"��✿���eh���D�YT���6�Q:����e�gŗ��b�\1��T��Y�G����zz����M��ػ~�q�{:�Y<���t�~&1s�.S�0��>P=Z�G٘���J���XL ����:�e��8WwC�"/~������o�
�)G���~� �T�{k�x��1	��R�	��� 3���6R.j����;�ޥ�F[�$��>YT��K�X�{8�\�5E/�����O��!���D�0�mW�R�8�b��w��.0����DO���;}�I�S1��ݘ\�\b<���ê#�V����?��ʆ�z[������pd_�ΟrF�+�O����P*�U�$1o�}v�i��:��0+��Z�3�;��׍B/��n2g2�������_�܉���2� ,�S5��dz���D@�^dTu��sN�	h5�4���Od��s�� א��\3$T2]�~�2d����$cCʺ{c��*�ʨ���w�aG�YRTX�a�x��Q�[2x�i=���ȫ�����$�O��(��2�|o�N�{y+	��$^��]ڝ�?s[<�(��#�ᬳ1�xUA3v�������K�
��թT�ꗒZ RD�n�]�Z�t�V".�R�.ȹ\��T����9�O1�=�k���@���!�
 �h^��ų:�f�A��i�]��F�V�Ǖ���W�]TY~Qhv~�볌�f4��K�&Rˮ?;t���ExYZ�j��b��K�
��Us�xN# ��顂e����'F4���6v�{��n^r��<�H�j����@ȴ'����Z?l\7�	��^s����M}�L��w������q���P$&��u��	|dL̅$gl������4�'�����^x�kW����i�i�����W�U$��Kkώ�MwMd���iD%E�4Pi6����kܳF��x�b���~�G�:�ŜJ��n��$bm�W+�\ؓx����y ��C�2'��k^�Ce]����%jwP�d蔍&ú������&�����PDJ�#�z��*�Z~�M�؎2hš)�j:�2�FC|�{͉�9��F-c@0>�shL(�կ#áK��T�Ɲ�R �w48�Yb|����O`��RRK�ifq�>Q��LӂLQ�A2�e������o�.��X�DIG����sT�]d͜/��������ߴ�C^#o�}u\�ً���h�9(�$ȏ�eX1_��Ϣ^Z���7V�O� q&R1��1`���!�ҥ��¾s9 �b���a��0
���V	i�&��-���C\B�|���}L�Ձ���Ŀ�������;k�,��V�J�wq��y�3�Yo[}XVt�;��u���R�۴U�;�/��'�^s�Ό�P��|��c�=�Q�����Rf����3���!�[^qD���5jJu��V�f�X�a��[2V�b)/w0��R�~Y�e��3�==�Av�wի�.}���,k�!z�5Dd�#�9p4�6u�
l�\D-c>eTC�J�d�I[	)/�9��)�VBi%��I=t-��|ؼ`vѰx���ɦjkH5��!*��l)�e��q9���?0N�����$~V�r��Ɩ�*� �+]X)瓉|���O�����M�ibl;���H���o|ya�cU��h�*��*��!�{��d��P�I��,��|S���_�|'���BH[ճ�"V�vCm�h���k���-:�N0m;�� ��f��+�PJ����f5d�L�1 D}T�H;�S'lOk0Qb�!F�vsd<�ѝ�ץ38w0�_�I�y'>3D���ο:2{n�V��)��?���x
���ADn�?�ߵ�a��L�]s�̕*MK��SY���lR\2]ssb��6,���*�7���;�j$}�%F�q͂���8iR����8Λ��`XE�D��E@�N"7bV��[�(|l�/ڀ%��#y��>:������3Hm��L5�5�a	$[Ց�D=vyg5�6�i�V��.#�w��4_�1�Q00�&N�{?ٽB`n|���%�U×L��A(}&�T��(�y���!dAoU��kD�7�&)��Mh��{eYÊ��a�>�����>1IC;Q�QL�Ƙ�q�/g�Xs�΂�����\��No���̘,�H�!��w�S$/�P���^�P~��
�����Fa"1d�N�J��h� sd c7�"�v|���4�ʨG[�;}�*�2
�8qNy��y�N���2����v�H|�J��~"z�X|�=W3��o���*ڴ#ˁ ���$|���͞��P�A�/�X�O�HcqT��E�c�H�8&gUR������=Ρ�����$�������QX��:�j5:�S��VJ�T<2c�Ԕ|5H���z$�9���:�������j�래eqi:x��K)mP�)9^H^Hެ`ڕmu��ٛ������Ցr�y�tK�3v��*LU�gN��#������v������z+>�Y�����G>ڃ��T�'�R����x���p����+�t#�� ����`�Kx�?k�=���N�ƍ��1,�����^��H�"���F ���e#�ʿ��>��š=����l��Mqlt�F���P^�ϻ4d��R��%���������_�([�)H��Έƙ�O��y�1W�L{�!��+���(h���a���c]Lx`Y����A�oyv���fy���)���h��,�Y�+(�v�27s_���T;"uA�G�;��C��km��_z[����8���6�3w+�X��s�=
}HTRc���|!���?�W]]\E'���@?�q蔀<q��<ӓeg^~���Ȓ;�5��2��//�~;���=���$�cף�B�hqpM���Y��骶��S��`D��+r�bh(�ƌ�aVtD3���g��#������]�<�ʖ��z��2�E�5=���)�XN3�&Hu������h�A]�A�A��dr�ө z.�m0�n�����5�o!�zœ?�τ#IF���k�����^��|
<ٳ�|_�WR��A�����w��N���}r��*�M��
⤍��=��v�V���K?hr�x#�|�Q�(��E/S9R�����c9���C|
`��!�w��;J6=�R#�{' ��sK'#'�����~*t���'󦼝�e� s�4�W�)V�sR�f�(��m7�n�\J�>.Έ9��KA3H+�1Ø��ji)��&�Xpy�� ?��~���Fʗtt�'zO\�
?�Кl	3�HC���JVv=�	��=x�ZJ�.��3�b�MV����EyS5�~D�l֎E��d�f�j����h��q%�rHO�&��������WR�Z�O�$A����_������DĪ@;������/7�o�h�nCP&����-�Z��Sa��lK�b��mu��ǁ�/u��#mb�<<T5|�%��U%���*_滟�Ǯ9��g����ie�Џ�(�׉u5���.A�%GH�n� S?&؁]���~[��儚������5:�xv���3,����وo��	���S�����1GS���(�Eg�ۆa?��2��=wzE^��*ջ�b�L�楠қ@w�k�zFJ�^�@k��&࿍	��cg�dD��^���Φ�(c��u\Tl��-�[��I�6(�y�Xt4�xi�RI� �	:cm<ͩ鮤i@ʮNz؏��]�ݰX��%*r��euwx�|3��;<ӊ0�!�.�o(J���n)���3�M�"`��];5{�tn���w�D���,LߞD_�_�[�=9Ž��-~`�Z%���ԪptYxט��s��J�7���B�`�@(�s�ܸ�;%��L �r�^	�;�:Z���M�'!~BXvx��ͼl�M��rj��>����Q�'@��t���x�] ��J
�7���3�xr�2m ����PIK�c$?�N2=�,���4X�w/