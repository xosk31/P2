XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���x[H]s����`"��x��,!�kbEU�
�t�4!W!�P;����C;Y B�ȵ���s�n���=�\e<j���eR�V]/(��.-��j�@&c��>IP���W�F~�y~�/e�~E;`���*7��,'��#��<�tk�_u��z?�^ǰq�9.~��lK<�u�#��O(�/y���s��>�o�,��/�Nu�E�;�$0NI�%3���: ]!D(�E�@u�V�s����eBB��P�{���B�� �P���m��nXD�q�z'jQR��+?TV�/5EƐ�?O�a��g�*!/�A�`�E F=%X�����#��e��p��䒈�Ř�Yx�5�>/{��l���CT:Å�2BUR��ah�tt>� ��v��{��!�p#a���샷Յ"#O�}s�@�!3R`��
�J4�H8��� NS=z{�T4�T\�M"7���p��Y�}�6�?{� �r]'  u����d�3�9��?�k��CcXԆ�4�S��`NJ�E��lj4���X��V��bK���S�KNλݚ�#Be�C����dwu���Qk���se��<`��1f�e}���D�2�GD�j����x��d���M��A����C[�@��l̐����6��/�� Y��4wbU�����\x��n�-�;Ʌ��e�X����j��lG�K�-BWۅ��:�;�7��Ԇ4��E]�H�O�%	�-���?)��x�Nœ#�<I��9�͝�G22�����Fths�XlxVHYEB    4a8c     ee0����4�h>]�cdk܆8���'����$#+h$���ؗ�:�
�K�p*7#wNd��nޞ<��!�O��-��G����`7�3�y%VSs��L;�:��-n��+���{����Z9x������pA�����r͗1�A�S_a���#g��#���>x��ye�O��=��sh���7�a%�����V�8���,jr��ò�}n��j����o�LO�_+�|��7�%�c���f��뫘���� ����P��������.���Z
+݄����E���:ߞ���f@�C[8�Ft�܈N�*d����W7�Dkٝ��b.��Mv����H�S�Au�����>X)0�r�B��kW�Mz���������|�/#s7���_x6YD��������Q�b��9����hH��:�QDg������ Kˌ���?��H�skFn����z&u����y���m'(`D���f�0`��$|E� �u��@@�3��"70���$��{YRCh��xz���!���HoI���#=
d��z��,M6[Q�$��-��J#w�N�Ҷ�P"nn���o�$��Z�*C�8��$� \�\|�Z�H�,t��!o	j{���ɠףN��h-�TAԳ
��Iʹ>H���ol�1`�LC/��4��N�)�͐n���?�Z�׎����~4�o�0m�����)�H"�#���m|�_2�=�/�BK��NH�.���^/yذ��4���n�w��R�Ru9����j<n���:ԫGO'��cˈ�9(wyw��\\�������~K ��##�krB�8�e�!��p��~w��������� {��0䁸k���#c\��j�w~������q���=o\��}��W`y<|�WgK�Xv!t.I�~_0\3@�ĺ�a�EC����jR*}��wE�HhDmRV i�Z|��:��ƪ�u֣haR���:`�1�y771)�p�(Eaw��|�%O��[�BǞ���A���.M��K��=W��s�7�t���FU!�j+�J4)8�Sg��P��>,VR�� ''��(U�E5 H���D&�"ː�a����tL�Y�4�����a�4���pZL��#ԕil��F�\��k���!��EyW�V�Y�����~�����O�4�`;��Y:��o�	F�Elh8��-����Κ Q-�IyP�7i��n��~����j0
�g΃'�[���-C���=8v�OUp��񕥸��hTAr�b?�A�P��f��I{�xF��"��S�D�7�hS��ij79&�z���4�� lH��:�O7�l�������\�Uh}�����Np��3�))�TTk�{�L7�y�D���+z���J0���Yۿ~r���Ͻ��Տ�-%&�	c/�}5ǥ5��-YC�VC�r� ұ��B�έ��j�l�/�O��u�R�Zѿ���eA�����OI�����_ԯ�CǾ:/GP����)�:�f�[���ۿg���%��w%�h.{�V������|����=?��h���uuV��PXg�PR�y�%�sS 2bf]BVlgv��X�&����6#>S�6�좉�y� ��:B����̻ߗ����Eуc�(P��C����PgH�Ww��j��[u����s��/{-�n	���<j[ћBC��#���&���.��p�^~Ќ[�0�%����8^�^�J��Λ*y��T6$#y��@�J��
��\�Ugo��rg����Zd���%�!Q�ƟH��{Y�x�}�eq��ӎ���Z�lJ���(���w�	��J-̲�Ko��)o��H�L�N��M�O*�2^.>rT�����\�bM��߳&������R�e�AP��9������ʡ���������'!�1۩�N��E��M�Zb��,�P����rx1}D[ޑ�p��=�{�����M�=#����(���qae��E��m�M���<�y#��� ��g"H�]�SE�?�������HT����n�kN]LG��\g�����Y������a�5����|�0�Q�� fy���Ї�X A��&&GK�rwYV��{b&S���|f>6♔�	)��X�N�M�	�+����7 V�GeVhqS��z1N	h!�hxe��`RE���cŶ4	�@2���@�:��:�R��� ��ZsMviC��]�
*����8��de��]#$��ͭW,�z���/M����a߉A��W�>uG�$<���JN���qZ^xB�8��n4ݻ��y�5��$��[�΁g��|���`c�z{��9H�.n-ď�s�d�oԏj2
�<f�58ІM�ӝx?Wv��嗥?���B
w-Z���I�Gi)aH�j5�i*XȃC{1z���f��_�q��� G��o�g��%�p���8����v(��=��y)L�
����Qӻ�+�����j�� F������z��G�Z���ժ���Fjo��у�+J������2�E���������7X���K�G�1#�G��`Ԑ�[�zz��#�}d�
��Z�H��g*j�]lk�Zg��(�}��λk��q����b����AW�c)A�������
h4Ҹ�0qt��	S8H+�hډ������Aq7�jq#�#�9Ծk�_ՀΉ�Ǯs���*��p��mm��5Bi�9���3l���.�b�$���5�79{��6���-|�a0�޶!>���i7&&}]�~� �xCg��h��EJ�[�#ɗ7U:Z ��ZX�|��i���*E�?�R�J��vm�j3,2��<00�&���m�����PL3E��	���5H�~&K鋇JbaEN����/5r��8�A�g+~�6��/ԃ�=�*`���+SV�	�yW����o��Y��8R����kK�+�P���s��_z�Fϖ���g��{qb+.�;Q9M��ûo?�6�U5����2CT�Ao>�<Ƥ2������n��7��.�R
�Q��,��O	|��^�!%wt�5-_
���3��M�}���}_"0�s�Z�+�c������S�S�;;�rJ�	�7�2�R��e�0���,(e��{���r@����\����Z/�X�[ �v5m���SXD�5�׾�<��0N�����(��b\��\Sv��mw��{3T��j0����
�9�� ˷����`Q�G������*2x>/��@�ʃ[%�����s�q���#�5H���sS��Wиu�Ҡ8g��"Rܤ��W +���o�2jr�	���H_:{����+U�!���\fxwr\�U��]�Qhf���X��7�qy�ۄ�Ò��HB��5����Ϲ�z	'���-Z�9��P�}O|���%*@ni�y�1"�p���ǼÕ�4n�]�Q��~���fd��V>����L�0áu��|{Ĭ%>/ �ߣ^A��F�c�I�m�v�)�#�x�`���$ZS�bp=|�|�&�K�~r=Ҵ@]�7b����]���vH��y�,ӿk��b����������K���$&V�Hd�����-����^������;�"`�1���]M�|�d�eF����9'TXo|!;g�C\ ���.)��ν�|���8���/�E��Q5�Ղ�1p���s��h�&~�2�G�N��(ˇ?�&ٷU����q�W�pZ�"[��%����CB�/P�JZ�����D0��O��