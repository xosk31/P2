XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����{z)��gd2M�r�-��3!�P�#�:X��{Xk
%���}/o��ȆN1�&1Y�"ر�u�[�[���t��/�y�^����EV,O<E��R�׽����*րf�S�|2�S� 2�?�(/��6�n6�1���\vα���6b ���?�e.�5%y����We1�IZ����f���J�h���	R#ܽkZ�@y��#�Z4zܩU?<�z��`�����"��tf�b��xo��7�,uo�8R��SfPr�����c�5�+�>A��\���.i� �)sz.M#����s�Q�6��i�Z��P3B�H�=��0�����Θ�NӼ�RC�b/8lJ����ư�0��Kel�2+��.!����,��,&����� �p$������0�a��]Dҡ[���,E��~����_�u.�o!�?�H܄�I��p$����4L�kQLd�I< :#�M��g���0��la0	��d<�*8��w��X��W���1��z�g��W����A�f�ω��Os0g�G�A�h4�R�>4��M�?|�V��?��g���FޣxL�'�%���i��zNxQ���E��b��3=q�,*iǜ���蔯�N���jm�H��΁���Y��k1����n�^W��3��[��N�Qr�n���GN��p�	�=�$�:ruW���4����������������Ͻ�O@�1P!�c�}��Y�BŁ\�\j?�Uj}k�����t�4XlxVHYEB    2f9f     c60�C熥n��}�y�W������(�r�v��L8v�sn.mX�v{�'0�7u�׳K��b��K���NO�v���҈`����rߔaڜ[��P����Ej�k�vl��TJ�T^�y�����2�>��J�R{���g���ZeKE{���0(hxG︼�����v�3��uI熬����4���������v������Ct�˶?2C��;�����Q�C����s���5�$�s֌K��<��%���D�]�r�3�:}*1fNY������L��uU%�^r{F���2���	a=��Ů}��خ>��X&
[ 2)��-�p����o͸�j��r���g�7Z�Af�V�Y��p#or�����D�;�i(��%
u�N \�L�p֬V��#ٔ�����d���	� r9r�32��nu��O;Ʈ�!�����fG��L��r�Ykr����(���u��~�ɣ�o­�&x��{[@+LES��Q���2��2��7jߞ��d���4��L!t>�61��[X(�ޡu#�V�"�a�Ο4e(<��>aa-�HG.�=;.�����g�l���j� �
���������6a��OF:�a�7�%�d��`�=J���53kM��,Z�����H�L�����Ec��A�����L҂l�~]����na�M��^r��1���É,�:*���2�z<�-H7Sյ�5kƜ��(�����`(���R �xۺ�����f�����+9�����R���Vb[H��<���X�`f6�ն�n��>E�-�Ϩ����(��N��������<V�\�,p#tO~T�G=]�
&��]�-���V�� ��D���ԴME�j+����D{� �:�PB3 ���|�b����P)tCHS��.��STt�a�����3/#-H[��rg�����A�g4�j2|8����x�?�퉞�u�1��ݐ�����q[�R��<Z�#gS��2|����d�o��7�.�x��j��cW�h�����˂�������p'�}k���qE?oC�)~i�π$5�I�7Qf[��)'XT��odP&�����yU��g0W����]���`�5	��s���v��%@���l�]�{�o]�J0n،8�V�,�<)�o���K���n3�4~��T�������\|L��* J���<#�2��vk��F�]�b$jj�_@>�iz��9}�W�b_� ��x�[�x�����P7���WŜ�$&*V?Ki|�f&����em���0 �H��l�|b{;�G����,�9���CRIE_I�.h��b�#0g��֢ljk��Tr�|�)m�����I�|�K�Torj�KH�H�b"G����0 ��چF�~�\P����-�I�d
���x6�-�Vj\v:H��7�A�"yjd\��.��m��ݔ�p~�oA�&� �S?a�P���t?C�+l�䋌q�+'��W����a<^�#����!��'~�.�RAݶ�������s��?!Z����ʚ�DC�~�O?�[�tA���"��Z�_�Y%I9/G/�Nܔz%7lP(��eo������+:EDC[<��%o�<�d�ޜ���  (!��Qu1	1�,Մ޺���<t�d�[͂>����X�0���V�7�=�䍹�<2�ө�ePi���M��lX���2�eV�f���~��9g�x<���K M�>@�У���n��.C�cb.���W�E��Z�q7��_c�%�a�-���zqn�M�xӋlA�����Ir���iD������x��z	�pբF}��}ysW�9�m_���hb������=W���������eR��\�P/�TqF�B��́��dzm�qy�9�����$5��Y㗵�ןeyɒ˼�tw���S_�$��Ϋ�	�o���R�������ȅ��m�t��f�g�"J���VQ�Wp�&-��v7��^��� ��U�}�0��������ܞN��ʮ��ka���w�'H��:3R��=�7�̨O��v�����O�`G�V"�t<�qs��}G����`E���P�pc8�ɳ��)af��1~)�;5[a��L7l��M��V�DX�	�q�e�^~*�c���.6��G\;Q�k�ie�8`�^����Y÷WF�VI�xZ����J���C���r'�a\�۔��|�'-�� �FM���-��9]L$��QhD��7G�%n50�n�Úg�1?s���i�#�C��ǈ�U\�
��o��#	��3GZ��	���@���y*b=CC�
4+0ߍ��d��� W8B����PyJ{���2�Ƚ`Ż� ��~~!�bv�Y�u܏��|G�4��mũ��N���V`ňag�P�����|Z�Ck��ð�:��Z�cn�g~��y��>۳}��hBf ��V��2np� Yy�5�5'�:��8Oo=vp��8eF�Oպ�T�Vv8Ryu��\y��"@Tx��y6����S�Nv�ɫ�7�vc��������z7{�_앫���PN���q�)ֱ!�^��iC��H �u^.U�6�>���ۍ&�zB�"2���T-���NV��@2�
�{&wb1�>�+���{��(z\�M�ޡ9����F*�KP(���wF������6��l��}�ި�PF�ˁt�S7��������B3�ԭ|rT+�Ny<}�}��W�|�C��f0��rr��Ǌ�v�z|O����tN>�?=����f�*���j�뇿��ӊ�ՉFj)��8�̊/W��T�nx��'HT�bԒF�&�j6w�GQ���J3�'�J%nY U�����F_�zt K[���PՁ\d���.{�#��3��؁!׷`�8 g�$�&Wk	�l�@��vi3*��\b*_��: ��GEK(���X�%����F"Q�Kl��l��hKAHi� �j��J�k�HN��3���'`��1a��3�� B�B�mYeŸ.�y�\k�ү={ȉ$��8�\�@��n2q��7�9�Ԫz�������O+����^���{2��7��]^"�"Aʽ��\�8��������a`G5�z���^��1>��D?�l�=Ɍ"JK���*G�v