XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��3��
I�������ۢ�vQC�Kz�4'���x  �<�5�����
�L 7�9G���H�E�(���5�U���zӇ���(`���Ì��V���yϴyDhޝ%����\T�c&�mG�̾,l��I�Cr���G�#��Y!��2ʓ��� >�ųB$z:���J��*?U�%$h�R=6�`Q2��*��N���(^�f$�Z$��jd�N���"�^஝��n>�HWT��i&#�8k	��8�T#�#H��Q�Մ+^�e�Ϸ�Q?UL�p����ݦ9�[�m�B?J���5��)�����7)r���C�WLo�8�}}R��w���ɁP 3����^㿡+�F;y����}�����!_6�G�c^�O�����~b���&%�Н�Yw�{/
�6�F��j"|���,lK���f�X�mÏ�0�D#�m7�<�*�[v��Fͯ�+^�c|��Nƶ�PZ�����psmxN��z�H&�>8ֆ�Ί��Pv�,����+��=v�?��ˁ����A�^J�@n����|]���0�h%@��bU��E`{�3n���f?���p��Fݟ����2-���sg�>��Pwiz�����Xc�d��,�gyt�~���<��h��4璿$8��g�2i��^Za�u�#��f����!�l�=��%<53_ի�����k(z��Z�E��#FͿ�1�"�"E.PͿ�<�QdW.�1�B��~�"X5�m{�f[E�~h�yP�6� �(D��T�SU�2��� <*�y� b2��XlxVHYEB    20a9     a60l��e��L��)����ˏ��4	�d���X8��Oj�W�Ҝ��2��/�;��Es��lf�qE�N���
�K�D��7\��T��h���|d��b�=y�5�_[�4�O3�_�"������o.2R�D��Hia���W]uP�����o�w*��?^��#�3���6��޵�dd�q��B$h�� �#P�����*���Ln�cdȋ_�(���M������Y�ﴎ48�w�TaBSgU�+(Wl�dZ�5����q���(#��f��~�#�n4ɕ��R�f���r;��B�)�9�%�2��w97/E��ä���;��S �����9��U�q��j�ڔ��<�9�0k3y4j ,j�̊2��iFi�m��h�愽��o��.�������X%A%r��\E���h�Jɬ9�U��%��`l�I/
z����>0V�y/zCp2Ҏd��[�z�t�Q�L�e;B���ds�ިM�u#o\n��pl
����,2z�1�s7'pCЃpH1��)��Ta�ѭ��F� ���9�y�g����^�p2�2�\^`�1����Mj����s��Đjs_���V��%.�qYܦރ��mT��F?���G�p+W�Q鲦�+����Ś�71���j#�bA��=k̔�
`�@�Uz}fO�����ڛ?m[N�c�6'��C"-t��go�!��5��܃����5/��1SS��)Z�*�����j:��;wɂ��裳v��n*Q�X~��=[e;��������Z����_M�}z�z�=;·z�������	h�D4C���:t�h��!����
j�4��*͇,qrra/o�uX�?�c�>ކ�hf��4��l�l4��|sg	���59�	E���;���_ +m�Ip�-낅	,�f�&
�Kl�S�gt��<Cr'׶�33��\����?���#�x9�<%��1��7"����`�8X�|��85c�����3Q�
�+�%K����Bj�GDa��l�$�^`��	�ӣJ>�p�VfS��I'�%j�%x��#A	���3=$�j�Za�(���#��KcC�C���m7u ?�H��֌����=ή|���{I�MhؐZ����Ue~����\̊#�ŋȘ���I�L�I��Y:޴�������lT΁�:_[C�:�h�h&�/���o���3��L�"�b�guc�)��#2z?5W����a�s��� >(�S��F΍��)I���{ R���<gL+K�i�.��/X�q\Z��i�ޛ{���?�CQ�z	��m���b
���NA��LR�*I�>���z!]�vC��?�iZ���b�Ow��CrT���9��o�N�m#� ��6煌a�Qw?����!aQS�?sX�O���O 4�v�y�11�ހ�+
n�j.BI}+������ x�J�g�V���N4�h�ޱ&'��w���7��2T��x�y�\�ӓ�-_�7w[�%��CJ�ָ�ꋃ�U~��Ey+����>�×U�e"-~3v:b8�z��a��i��*���M6xX7,��hĳj��j>Hq�"q-1^\��M!�� 6�ɼ��D(�`�-�l��/�Q,�"�䜧���E�
��F�	M�#\r
��]bP�S8v^o�Uq�Gl���̊�M�?�����7p���~�>���������#�I��ə����"��:��琄\%��$��ۡ�Znt�@x&ⱡ~�.�KI��޽%Q	N��o�Ej���\�]�����,e���%.	/�ȣ���X���
mU�~GA1�Ƹ@f�0
����ǩ�~��ˎa��zw�Ze��W h\��hUM�D<��|Pm؋��b��ր��!r��e�h���O���V�X���/�>Ť�P}'!p�C����X��K�f�q�V��O�+�Or�l�?�ed2�O^:J�|x�O���-D���c2f0��W�黬w����`��/��;�83L]�$k��bƮA��t�O�b@��rv�3A�jǗSq_яO�&^�;'�3��X^��f��\�8̥�@��\Jy�኿o�lz�O
�.?t�1�Xt����9���!6�;����)�G�
�_����3�)������p4��p��j�����
�ՑYUi��5$�l�W��q,��������e�N�Q�J��}��]n� �;j(X�2�T��b�M~N2�bNч�"��g+��ޣ��4�����	́tGR�}B�u?���|` ם��3qc�ƫ�h��O䋛������>4�_(j2�r%s�,���F�w�иZ1�ayX�{��.�q�ʜ��#j��[{�r򳑎R�T!�w��Y��G� #�;�Zݾ�|��DC�q���}�I���/�-42q��S��/�k�;E��\�$�^���_v"R� ���I�zg��7�r��yT�V��.kY@�ٶ�o��#s��ª3~@$ɂ�����s��>�h���ڦC�y���=B�%�]��\��	�c��Y�WMpD��4|6�����V�P����s�O����S���͹nq]-5*�Y�K����K��a��B��Z��❌fg�w�|`�T����	x�΃��t��B�ac�ES}l/Ed懣H.�