XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���� �Yʛ���[	�6���{������ 
x������<�]D�x+�S8������ �jk���Tk��*7�b��'���H�tz'tƧ�3<(�2��LE�9E�U�5E�q5D�H�Y1�s%�bC�{7)\��`�z�D�|q�;�B�Ss��q�y��՞�Bnlk�}b6�ƥ�R� c` ��w��i��m��͡�₞�k��Y~v	��S����Xb	��Ң q��}3�'#� qu�M�EF�S<;S��9�[v�[�ÉO�tfv�-�:��\M�ʞ��� �?�(w\>���>V�����y�H�[������B'.�U4_#/M@�#�R�а2��$��A-
�L#:
�n��^�9~	a�a������-��S��L�D�{�<��dQ�ǥu>	v3��a��
Y�?��W��;�1���SY�Wj���_1R�0�����
a�Q<A���}-2�����.�����I�N�,8�SEP�*��$5^���s��|��;���i&%�)�Ǜ&]�c:�z��r����VO��2̟��gO�����Z�7������8�ǟK\��ܖ��UM�}^ə�q�T��:��3"s� �DP�hG�G���աdU�b����Dm�������*�9)�biYף�?��{ę3z%<��W���0aj
=aR���rnfZ44cڧ_�f8R�o>�t��	Ox�����k�d`��P`q�d0��%6���˫�� �hD������n��;�u �XlxVHYEB    4a7d    1090���/��蒌����ȕ���%��v`�t�u��{{���}��ֵ_3�`�^ʋ洢����{}��F��N�ה ;����d�;V�;�ܟU�RU��!�����Pc��_o���p���q8QfEtncm*˳}`��.`�rP��?�m�j1�'V^�^r�f��������G!#��
Ӛ^u�Ӏ��s6�M��ϥÍB�'x�i
�^'�JsǤ.�]�ݻZb�o�:ZL�c�'��G���II&JG��Y��y�=�asJ�b��?p�~���I�K�,��[�Oz�ϧ�nC=��O�зKJ٢�ӓ]��W$�7d)V�Z���d
�P�\�a8ܘN_���x�^ǔ��_qN�D5,+�'���d	�{�1 "��Y�f�ED��N��q�ҡdWĮ�e'h��U7��+پ��{Y��PA��h5\��`�Tk>���ֵ�-zkg��H|�#9��C.N���6o9���~uJ����Sc��x5|�TJ�ٌ՝�}U�U9�کC����-&��)�L��|�J��p<��'D�����Ě�Ԛ8��k�Zd2�M�8�gՃ-��H.C��7�{��+�I*Rb�%QQ3-�2���᪃'ǲ����%�o��Y���<�2� �x�pc�Ə<���ŭ�qx��?JW�g�J��7<b˕�P
~t�e�j�ԣ ||[���j���r�h))���Ռx2�	�����a+,�i*u�*铼��N��P�8#�r�;�9�<!I>L�����`�*2}��g��%a����W�v�-���mɲnwE��a.�s`����d�?�+�/A,��y�X��&���'ʄW�<Hj���,�w�A.p��~��ֈ$?[x��jA1�m��5x�6��'tTD�xy�[sؚb��,���x�,�Ly'p�a�|�?���PN��e"B$WT!L	)�ޘQ�9��8��ڌx�}�VOx_�bf��3l��IjI�9�~��M����:���HG�O��:�6F��4Q��ܤ8�Y��c�k&���R��pO�0k��o�G{��;�I���4�gj��40^Qr[+s�1��L)
�R������N�����d�c��\ԫ�s�ú~/��=�����4�l�<�ۑ�#�M��b�Bg_�)�{��!�)�+V:�?���:�QVEՒG�������5����6_B���bO9�V����n��Z��z*�4j�΅\. j|7��uT��(�t~�+�b�K#��-���`g:-4�GZ�ԮG�[��\�P�{ٲ*58�p�RY��q~K�C��?���4�V}��і�ԦY"p[R𳌊�"3���DJ5?W<Rq�YH!x���v���[�+�Y��#�W����Y_eI���=��ʛ��Υ�{kASm�@��k��h����(@�B�awBN�2��R��@_�w�1E1��z��_�!%���K�d���8.�H�S��|�D���w�����]l����?j�@�VX��۾��w�Z�;VV
0b�
��@�8��~}�h�G9:��a�Xڽ��p�6(j��;��ϕ�HNGn!T5`Y�f�"-࣪rc��'�U�J�����-_�U����ah#<��N�]P*�\��U��o��Z��T��l�#��E�³�X�3�L��qזQ�}��R��8� �^�AU3�İӷ� ���L��ծ_9T���ݓ�%�I�lo"˯�x4�;��d'�q�c��}��n�����F85B��t� ���]����@��0� J�|x�?8,����08l1�x"��M�/��mQuB]�q�,��.S�ֱ�y�Q��E#ZCR8P����I�Ȍ:��ǎ�*�#߿]�7yғ��?�M�g�ʪ{��lꔂ��T(*U�qmq��+%�K���i���Z����c�$u�E"CY-M�%K^��m�t0fa<�!���0��N�#DViH�e�8��q���ۑ����4.�^G��x��:�W2U2h륿��"�،�ԋ,ɨ�|���w�F,6L���-ՆYX�'9ӫG�:��O�ۣ�j� ���d�q�m�X���/�U`�҉�}}��(�Ոw�Wsv�#f
Ve;5-|/u���wEA�\|�lN/ukE��j�P�4b	�����d�L���(Υ)oi�\=;�w���ZV��b�3�b^t�Feö/%�����
�3�ٞ&1�>�q��-d�h��.33�y�C�5�S����vL�,y�a��`�#�� [�����2c�p�b�Y>����X����ӝ�ä���3{�s�mE��O+�S���B�E��@����C����@��|B�������k�1�nC۷~��'׸ ������Q���VC.	zt�v,?��a�������>��(�S�5�KOT�z�P�௓c�^�.��D�wAZ4�p�5b6������H
$K�$(I���tF�O����lq��ZxD껼��}����%VQ��Ȅ��U�Z�L3E͡���)�
K�`�#�*���������@�BT��q^���T�`�HLU�Cb�5��I��~�~����q�Feۂ��(y��A	�ʫ)[a)�a��=��ە
����*��`��l5������ǒ(�e�h�g��;� �3�<����~��'l|���>5��>�WZ��h��I���y;ih�_p*�\�!��g^�vw��K����w�3��G'
�P����͕n�2(1A�H���lV��L(L-L��/�P���)1�/|1����<�vR��V�����p����V[X�N��k`�lc1��H�a·�����!@H��בc�?�D��ԯ��
�ٰ�)c�0��q��$`����A=�}�����8��y�0uL�&�=N�*�$f�L z���<f�+!�����#������6X��r�Eʿ�|��0#S��!�G~+4�َ�i��m�����}��$o,+���D���`:��/�t�gL0D�������o�,��=$��t��/��7�X���m7��$7y��Ch��kt����PF�:�������(��E*�Q,��j�b�8�<��,]�!t��ô���E�0�͡�(�m��"���ۈD�#Z��OR}VD��'�pv�tԠH?oY�Y� q���i�5쭸�u��[��J�x�o�=3�1�� ���z�x���}E���%��e=bR�PÇ&��RP��69c~�981��Eg�3Q���>I��/`ŊzJm#��h�|Џ4.y���hܽ1��<�9|ܧ��q�<�!0�~ⷋp�Fg����Rt���r��ͩ��i�PE9�m8�d-5t���5߼hHDqA$Y��*��5_��A��>���\L֊��j�ѽ�4��XU�GT���3E�L�s%�7D�t]zn��R�)�z��$�I�ZV�qC�z^�ۄ��0vH�m�R��'&#5d�L����{�R	�^=.�-0�Px�S*��8	�����{���@���[����\��̏�A�5�l�?a�gmw�Go�A6ܮ�-�-z�������ޫm�`��p2
|b��O�Z���m
A�Tː�������`��w�B��K"��d'�0�$��Ҍ?�����ϑՉt�����U�+�`�)i�H*>Y�P�8WS�WJ�@�S6 jm���H�S������\kx^�RN����s�SI�l��>q�Jx����B;���nK��|�0+o���:�˓bE�.G���0S43�׵DM�����(���m�h%�s����+��o�:�݃����>���'?����twVv!Ǒ���t�(B�%|4N %.3�}ͻ�pfP��7�>���)�S��Ʉ�ː����f�pP�j�7琀�ȕTn�F	�:V�cJ?H�+cD��G��w���d���r[��1Ü�+E��s��c���Þ���W�&^��y%�dKFt"a^��t�ⲧ�'6z �V�1�oV����$�e�.vQ(^���ؓ�\+��M�~K	����
On+�W�kE��킎�tx����}Ѯ?�ZBu/EH���d��s{4�am@3)�o�v��ylOŔ�����YS(i]�Cm�-�����3���r#G�sH4Q��11�4�7�0�Psk^N[6�������l�/c3G�a֔��%%-s��!S�����{i1�]Up���Wk"V��J�&��