XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��RZb��=A�F�
-=-:�����%wH*'�E�À���'��xû�?nW����u�p��I���{�a��m	{��ƥ~���]6f��,y����ˬ֓8��M��R{�K�+Y�e�)�w�2S�%�lS%�B�3�+�=���S
C������W̏��ݸ����-�}@�'E�K�4��?�q���ɅݯAdv(�Y��MG`��7����?{����� �(�f����
b������b]��m3�,����ĚMX�A�\ް`�I�S��v�4.P�ȝ�R���;ƌY�$��Q�٩�zc[�I�V] �]*�,h#�]�)�o��q��l�8���ss�q��mqx'��G{n�m�_�����8�؅:���-́?�繀'���̲+�������<�̗��H��3�6�����S<8͕�LOh����\���ӿV�N�ms����hz��,��3rUy$��F�l#Q�M�xE^P���A���G��o�b"Y�g�dG���a���NyL5��f����=��߾�Q�zC����ٖ�i��D�]K�̈́��-�/���:<ٶ����s�g�d�6��b1��E`��]Щ�`�I0��V�@�}��7��6W@B|���Ec��؂��+j�6#(�A�Zh(�ER�\�ngM�B�2����C���>M*�!�	��&f"a�>ڊĄ;�㺍e�;�Q��aץ�,N�]m�	�����޶���٧�;���>,_�Қ�YP� ���9�bt�XlxVHYEB    549f    1060�[^l��5���{���E�:�e����wdC|��w��aKad8���@�����N��Zm���bx�?Up�{gS�hop
y�����~��*�SKo_?�H��iJU�����F���I�������¹�/�>���sCթ	8��i��G��/�>�X!�~�������f
p���e|�	����B���nD�S3KV��v�g`�d􎮍s���Ȳ�x��+��EﮧQ:��$��Ϻ��vƐ]�/i�dx5�O��Uj�R�
f]m�R�bxD�])�Y�ͮ(T�c$΍�w�
�z=hw���R��Ctaϩb��Z��0�_Dli�/���t�j&D�]!ʨK$f�U��L{![�l�L�����z��j�u�l�L��~�����"��a0�A�;9Gxz+�/l����?U�H��o���8�^��v�y�E�u��P䱜h�w��YC�_o��,�S� ��"c�G�a`��p�>[����/D���L�ڱOǇ5 �� ���%6�!�����bi��I֖/6�&yC��K�?v0l+)�h`���:�E�2v�YTX�[)���5e�F��Y�JL�"F�5K�G���ǡy~T?eu���[T�Ѷ��N�ߘ͢Z�=\t��0��}a)�������L#�|6�E�=�ׯt�����~��Xu�b10���JJ3��:D�(�8����7~���{��X�|����F?�(V}���6o=��^����[h�PۓxN�l�r��򾛼�K�J}�#DK�"#?*sb	o�]X|���'��/d|���5����<��$G����L��A3�q����5���;󼰦��M'S�ȫ���F��M��B�UCS���%!��/W��8��|�ٙ�&�e0��L�mr�����cbx��gT��>�!���w�����G�>m�p }�Cr�^����B�n&�@2K�7��G\�2�Sl��)%r'>�N�|k�M���76s�f���	|�>HX�	�?p��EZC�G�Y��ܳҥp������e�"*Zݣn+� ��'�������&�,&��z�{XD���ͣ}�y�7�_�t��-��DE8�(��-��T��"ɡ	�a�1� �X�3���	Ҕ垟ʡ���E?d�/��P���8_�=]�
���v�ej���&.�VS T�A"��R 1�0]��S�uf[�L,��H�@l�I@ 7I�F����	�d�A��҇���QF[iA�Q*�0j�h���@�l��(���M���nk�X�w�[z�������L�~�̻���f���+~&:m�]N@���/s�%���$U�P���ϗ�U��[�!\wEjש�lY�)���o�$%��=��;OS|�%��� *pj*�g�ˁ�������p���h�9���ʍ�ՇK;�qYrE�k��N�<�DjU�>OќypXW%l�U�k��<���D=��R{7t�z���p������u4�L�����"��H�}�]�^3�� �5|�k�6ҹ��C���s�[�&e�Q�܂�/�<�˼�_~B���0u�ζ0*��i}OٵHV�
�����wG��PZ��a��k1Ӎ�v~yp�*���2����YXg�Q�Nr����t����T�/߅@"�Y��d���R,k/��]�O�X��h�q
�:���"@V�<u�s,� ;��w�r�:�s��v��IyQ)'����'��OA�/�he#���$|<(�o˦7�<���u���cS�D����D�j�z�Hǻ�V��ӭ%��'��M<�Gu�.�S�R[��Q�X���!�*m�\W�KT*��Y�H�F���q��֟Wzp�|.��3U~v��"SL�ք��� �^�	��'`���B*U�r�N�<fPJ�a��b6[�����ň~�(O�)�Z������#�C���\�|x=�&x�]�8�u�E��A��%�^K�ɇDlعe�̽�#Ss~iW�0d�=�V�u�^����R!/bX����	����p�VS�O%��`�W�N��q�|�꥚ƙvu%@��N���U4�	�=����K�YW�m�$�^ƙ�X��o���9��Y���P�0Oy�Ո�e#��ZsӮ��v
���O�%���O0F�{;
�-	���-��7���_c(8r����(7~�������S)Y6N�?�ҸLǱ�����'l�_�0}VP�'J%�R%�<\$���Д�F���`,�i~��=3z�޽���pW�=
���.+�(x���/�8����e� �w�ck-��V9=(�o�
��}�v�i-��f���O��q�IaG%� �O���Boœc�.t�gf��lJ��dC����Fo�ZZ�T��d}�NH��0���.%3gͺ%9�o�0,:��JJ	�7��<����e`���K_��`f���T�>z���{�X�	Z% �JF�L���V#���R"B��1�� oPN����X�g���n�Կb��;Fr��`��ce�-�����)c6��K�6�U?3pa��@&E�*D1Hg��vC�!�����T�H(���8��� �0�'m�=��J<*����CY���2��G�Y5m4�B|�E��b2�0f`;�~��k�,3��ފX��1�h0����Z4#��P:�9673V{�B^��������.��M��pD��Y2�g�5��PALQR�74^r ��hy�A2��:�j��f���s��pTO#�
�:H*r�O��c�М�.ݓ�a��V�O/�����	�n��6(�6I�Zh(�8ҸC��ɕ��I>��l������L��y
U���]4֒]a{!`p��ܵ
��v�����e
7Y|ka&��A�<zWÌ���sc�pF�j��r,��7Y�0��_�e.Ǎ��QQѦM��h~��szՑ�������e4�
-�d�q��S�ᬰ3L��/@N�3
yފ�/�Dj�#b,��j���l����RX���3Oܰ�/L׽!ksі�Z��<��6t���1p�Rn�X�T3�h�?����Fb�WE1R���Z76��q	�Y��.Gs��3cp��٥�dGc�<%�c����-#�Dd���,A��[C��ڵ�y�w4%��9;�Y�"�W� ��������h��z����a��4�[�V��S�|B�O)��0����QG!��sx��le�huBw��c>Zv><|�x\��~-�0S:���P������S���Q���	N>�޳�9���OZF�=��c���uǚlNs[��&����Y�6��/4�,k�E�re5�Xχ�+lyuŪ$���g��t���[�3Yd�����d���C��Ey�v@���>�lq�_��5�~E Y6��I��<DD��LA�G@�v�73Tȃ�� 3�?#��Z���^o=�K��ֱP��y!{�6*��d���	�9��5�"S�&��E)��pEK������b1�~EfA��e���gܯ�!=ԯ�5���yV�k�`nj��#�>�[��t=�vx<�j���2�|vo�3rE�)�JQJ��l�q�p�İ������\�E?�ګ��mi$��l��Ԫl�a��(3M�8�O,���?��^�kd.g��/
4f>̠�(v������bL	r'�*�������־�J�62�&�bٝ�9`O�=M�/�D������� �rD�C�(=bM���g�}r:�k�
�Λ�O�����`��C��	�D%a/FS������R]��ļ=p4���:���<'�A�?��{L��`u���R�p�)7`Yn7xcS�Xu�ڮv�^�E\����#�ƴ�RkQh�p)]o�79�\8D]4=WwHmL�$�Hj"';� խ*���ő��h�Q�bڋ������i�FW76S�Y�P6������Z����A2��:`�~H��S,r�C"�D���5%�+jx^6	
�8�l�6�Ԓ+��}�>�H���mI�*X;�e���v���=Bg�PP�6@�W�}�k��*������4o��nC]l�X��`��ǵ�|'�*����JAf9��גOB��Qap��N�H�0���r�p< �,��Jd0�x� K���+� �F�5�_3SC��HAa�l �ڭ`��**���m