XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��@��D[��Qn!b��m?Ҭ���u�,���a��Q_/E�r��%`CGM.�P!9�ݝ�����8ަ�+s�|�עcn��~]�6�0�������j��G�V���,�`����%��2�ſ^*��r]"�L�[p�iJ5�A�?�Մ���7L�wwۧ�t֬�eY�יq��oj= �?P9��9�Ű� M�#bOhQJ�Fݺ'���h��55��H�W'�48�a@��0�v=���,4�7��zu���_��6��Gҋ�lO#m��R� ���Sb!:2o�RO'�%�;���%5�¶Ob}�L@�����`������#'�k�g�u�Le��;Q�qU�#�Uo����̃p�ލ�\8IA�0��+{GhsM���˱Y@3=���&P,(r�J����e7�k�~xb��N|I��k�y���UW>�����r�ǆ�j���Uz�땆éF��g-vV�s�7:\�n�uE��0;�)�<{6�i��v����<�+�[J��ڰ��%+|�
ogû�2a�e��]
��L�=E��FC���i���G�c��v�(L� �5T8ßy��a�x�.����/�o�WsX���������U�-w�l_�w�s�co���aw��e|����="#��C��Tͼ���;[HIy����N��H~}y�I�`�wj��-GvǬu��2�]^K��'5�k��`0 m��W��,�*�^d`Ɣ{�ڽ���-�
v���2��}��5=ޛ&�e>��_B01���XlxVHYEB    b8a6    1ac06��|w{�6�o@;�H�!Hymzw-��y�N��'�6��:�P�0R���U��4�X5�k(���3j 5����*��P��)DQ���iJ�m�7��)]���kP��:�*���h%:g��e�ukە����5�)A�͹�S��M�\>*�w�Z�:���>��R������h�����M�ϙ�,�G�pk߭5��/o���e\��v.(���h�k���P^�0K��JC`Qt������YNI��@[U'��·:�.��2OqM'�jC�9׋�.��&�ɺ����Cl��g���!�	��l�(4���U�y�gM�۞�)~ L<��O/v�k��8�8�P���
gՎ5:�Y������o����d�pJ��o�f����4�ܜK�^�7n��_}
��%���!B����R�N1�7�I�[�2�fz�F�zT��6���"�����[gط�Ƌg���_��s�Y`�;�BX��{�Z饑����Q�S��F�ш����v'�]#��j�)擪���Y�;���6����^"n�r}=�Ff�R�T�tb�Ŏg����H�J3�+�B�����p�:����l����	8�3�b>:��4�ΏCh]�t��枉rZ�*9�J�Yk	f�,������b=kwEj�Z��U��f/p����JIVq���r���F��.~�NU��*�4>[�nz�SQ':���Km�#�~5�H��s?{|Y��Aj�������G����J�O�-��(`������z�hh[��כ��̏8�**�SԲ�K�ч�CQt�� �����y#�#Z�a�`�k���M��:520�^�K��9��LԸ�6�h��^e�m�U��6��%Ȗ�P�ۢt�/��f�+���I���d*vF���<SD	�bݩ�Npq2Ҕ�ˍ-quq�Wq�9Б:�����y:�!�>�j��iy)QKoe� �]>%�o:7��#�F+%��V��V��5����~�* �~-)�P�A�'�H�Es�&��(��.��*�01F'O�Q!T���þ������mؗ���8-��-���UG�������QC�^�v�p�� !>�z7+�_��bܻ&���I�D�{u7��4���<����#��*�G������U�8E�l:k��=vhl�����lD�A�*���L���zu�d@=*��}���A�5�8�PZ����".��_e['�{�{�iOu��X�������;4�"+�(]����VB�K�{S�J��S� ��H�ԟ~͔:��y�'�Z/-s(]��)��.�?��ћ0��2'�;�5�&�;�Z�cA�A��!��MZYKb��@�Y�w,F`�4��gIf@�x�hU!<$����~�sı��:���x��q\�?���F%�#}'��*^��[P#{ՓK�.�:�"Ԟ�^���CiN1�!Z�6)|C6X��l�@�B�7��s��帊$+�Q��%�e���c���8X��Yj�d����gl�[�GG]s�ݓ��7��#)za���}#�v���<�t��sQAx�c��i(�і	���vU|������C���;�w^ጃe���y��R�W��H[۟Л��c����ƃ+x���uI�h����@kw�dh���>#"��
xf��nA%�	�rc�Vm��l8�U�Vj��D���Ŗ�N}��&0^^@���V$�.���s�Ӑ]?%��~��2򜬀����X	���Hu��b������/�L���g.D0j��1:��岏w��g����`N{�4U�8|xF6h���g�7r�6bkr��_yEs���r��?�"���ȺlYʯ�-����	A�	�=Y"�\���Cՠ�o7�S�Y ���� iez"�!����
�t|���+>j:�*^�MZ�)\����_Y�.�Lfy�����j�>7EwH�����m��M; ���|sB%m�t
O�Z��f�NX�JH�3��pIv@�H�����Z��_	��s�K,��R���|��r�n4�(@�`�4�#Z��xL8�Q�J��ׇ������t��a�����\�-��F����L�#(I��U�dI��F���%c>ᔽ�)g�o�/7t��Q�Q�*T\d��ڶ�c�d�b�n��ZӫG�9��b�ٺz���ї�*�v�1{�5_��(,>M�����O5�2ga�Z�=�\��ɶcf���<����T*�L�٨5�?�����?���e��>��h�J�v} ޿"��Uɕ�R	&ܚ R�4�r/�c3��m���OB�7��
:�&�����qil��=F*ѯh"S�Y�����]ԐT.��"�x3���F��\j�5�p�T3}�&����ٶK�%�*�O�l�#��{�\! %J�7���<��`�:9�+"�7��n�����7����a`�	a��>�6pì��W�"�>]q���w-�C�k���'
�h�$tn�O�I�qΑ�(�I������)��=C`e���ŗBoں�������!E����/qg��r��$�G?!�U
9����I��'�_�Ѥx�PRk���c�
� 5�ȃ�)�{2���r���&)o�0ƞ�נr��8��^"J?/�eR���s!�ㆅQ׹�,3��`M?dЉ�q�zzP�80��ȋ*�����gJ��9ڿl����#�ݛ���h���?^HO5��_X=B�����V����E�A�S�G9���b^�������v"u�mud�p�#�<H�᧴���eݞ	R��Eg�_	k�}%ɡ�LX��F�k�xO���%��z�c��*\MA����
��Y��;�c�����{�%���$!�x}�wmˈl�����\O���[L-�bB.w�)V�o�f���#�bdBC���*�'u�]��;�q�Y���ЙZ	��2���o���)#c�9��}���;��G3���m�oGT��v`��(g�-!���~���c[������sX:А�ʶ�8�&Xگ�Y6��j�i�	��j�E���^�hjA�(cO�ޢ>�bO(Z�Q�H�ox��u��.���e��(9���O|����T4I �8ʽv,!׹
�x�T
k2��-wtx/��ye��=b�UO��j٠����	xd:�H����S;ox�,��l��27���4<�_�<�?j:���%:��x苒	�"�|%*N��FG�Uv�]����x���AR|6śn�#:�v�X�p����g�6�G��bG��K��Jgr�|��zO�R���ZE�4�E���/m��[�_0?[��j���x��|��ో&X�Z4�'�t��W\������_qC3�S��O^.�6�� �V}�dlь}���~���lO��T�!z�x�Q�hF���ڠX�b��KE;�!}�۲$TN�;��s�5t�m8��ګ62~r΀��t�T�;�9жv��,��Τ�A��Z��&?��Շa�S��wfA�58�|( �%�z��6�N�ntX�e�;틢�2hyp�Q����y]�Cy������B����q Beڦ��?IBe�wL0��6c=������6R�%= ���1�C�Y���p���rxI��Ox��-���x�B��"F�W��a�	�`��$�� ��WB����t/�4m\�Iq�:�v������fZ�͒��+׽,���2��Q��$3:|�&�:��CN`|��^���Iq��i�\CJ�VC�`�]��l���~��Ч����(ys��S/���,+g��5ڰY%�4X����|���p���������&g�Ӳ4���h� � ����jS�x�X�E����K$ݠ�0��N��/2���<�B)D�R��*�eF��\@ȴy�	��Hb���l�V�b�g:Q�^������d����4�:Ge�� ��kQ��P���y�Z&N��؜|�#�{ ����j�+�p�����ż!Fk��A	 \ p��<��-�����.�w��Rߧ`g�*��Z�gw��H��{�/�㤒0����B��J.o,�P����Kq�UtH÷�hG )ɹ(W |sy��G��T�\[.�m�V&�K�~���Ԥ���K��<�*l�,����!Pz��1k�E�%)w��{���p��Y��E�ʡ�C�~�Kۃ���f~����6��ߨ۴��S�ҙH����o���a��m���&ޟ��\:�`��P�Y�	�L*vt7����=ˉ�X�h;����G�,in�Oq*�| Π�<B�`n��G*c�����PV����47u+���pDsr���G�b2���7��B�L�L�Vp�hI�u���|\�9t�����'��Ƒ�Q�@�b�����ֳv����q��uu��N��1>���6H�et�a������"X�c�>Ag�&�~�V`!�4�����;���/�Ԩ��\�j��e`y��@H>��z>�&���MB�y^�z���r�� ?�Q�7�ܘ��\��H)uDg��w��їg�B�����"؅�*��F.�!琂�)���m�F��0��N�9NK+�py��;}<�q8*N��L�r���΢��e�dA^X���+��XA�L����C��xqN���t9�౸��<�.�c��P���ɉgfb��A�lM+�ڣ�	���&�� �����jK�P�\čio7��E�y�>f������4��4v�.Ⱥ���`W�.��,�loP����A���4�M3z	��߄i&�4�r����p��QYh����p��*6�#�`bN�Sm�8��c����C�����cig>_�s���_��&H�j�˱*��Y�ws��撃p��ǵ{B����������q�^�F���RK�A�#��9A{�!q�8���nN�[�
���p�s�Ǎ�:,U��4ұ۸���y}l��2!k�~���je�2a��M�������-����3� ЀE��$mt�X_�/�)�u��+]DVYc�/ ������[�:�;��D���C�p�GX?�f����!7\���#|�����Վ|���@�$��.-`b'���7��(%Xkߵ	>��f({AYPX� �9��A1�Box��p9�7�48qc�3��Tk�el��E^��5M���!�^: �-%5	�O<���̥z�ރC�;�4|������2���l��ku ��'�A��=x?���*����WMJ5ar�Z
ɉ�7����̯�8��H`0���-Ӳh��B}I��Z��� �n�`��5>OGM��*��9���8&y�ꖣ��*,�p���[��r��z�9&e��������b��Әl�a�8���:�n(�Z}��p&9s��6�[��t����
���h��RG�9'�"25?6����|茽��O���I�`��ތcW��{�Nz*L.��#O0Tny�Տ��?���;_��Z��Eö�˻���`��W�}��=>E̺0�Vfm)�-� ��W�\���u�P���T�1쵬�
���rC���0�lj�Ȯ��n2���5r��J�ſ��;�Í9J�ӯz��Gɗ�p8��#����M��n��~��P�\�J�>�xp{�kǧ���s[��(R�B�GZ`]�^�D*�]-?�	|v�9��[�ᬧ4���8�YH^��ot�_Ս��dpB՟s¥Ro��`��Cdar���6\B����H=g'0M�������q����iE��>Rf.Q8H�}EX Q�@�wQc�~:�dHt�x��]-�^���(�p��;B�yT�."�o����������KG,�F�0����'+	����8��V�K#����$"	�4�(D�U&h��$S=�G��ړ�J��Є��_�e0��S�N�2����4F��s�I-�Q��C#�k�K���@�����vwș{��4)�{����9S����^3�/�0u[F�����v�EA�Mϣs�nE��JN5���X�n_���5��ǀ?̉�,��B�U"��Y3Iv���O��:}��XU��Va
�rZ�eXo�ƍ������"~�q`�j���ӗ`��)�:�� ��j:Т��+�}�(�=p�6��;��Y�)
��}ݓw�!Y�2�$�|���FέԺ̣F��n��Tv��5eV�&�'�Ox��؋3J��Ѻ��Ǎ�^)���A���+��03<~7��_��u�zK�C���󑆕�������L���5�W0�pU��	���n����$}�]���2����������E�+f���~��v�CgՅo7��h�9�(2�`�#~��Ҫ�$�43@���$$���K)C�LP̹H�ǲ��:3e�g�����'�*�)��_[���Y�6�}F�ȤA�u��rX55J�K��ʉP�w�1��/ ��9��������=�Ɉ���I����hl��.�$��0�lE�Sm�� D��z�}���ޥ��Y��'�*��� �963Q��?/k[�{:" �ޏc`��0g � �J�cݠY<G�u5����e�i�V"��A���m�/�B�/Jֻ �q���q�"��y�:l���:�J�
_���S��e�i.�ȃ���|i�Σ.���L6,o�G�f(�Pi�AY������)G��E�ͺ�M���BC��t�;X`�65�rr(�>���dsIf�2���Y��FN��>*'c���M؎f]\����{���$��PHYN�%*��G�1���1ǵ�m�l�W��gӽ��V���6]���y�������D��_�%M���3�