XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Tg��V&p�@�c�#��*�j4>_��W���`��fQ��LK�)�Y���<�h5\�w{t��I�����b�[pru]�M�9/�!���^M�V��� �T�2�F��)#t���ۋ��gXj��#`�"��=�@��]�4"� `1w�Kf�ŚIw����kc��i~�L=�>��$;ʌZ�)ʳ0��U�PX-����$F����ú��<s0Z���R;��X�V�����W��P]Xv#��ܳWKE�Y���d;IW�ykx0���	��Օu+'�B�`ij�|�8g�c��)�h���@�w(���H%�V�hb�t��'ϕ90���#Y����U�+R�6I�w����&{,���S�^���;m�d$!���84 ��\�ï�bE�W�p��?�{�$OЃ��qD�ٌ���$г7����m�b7C6'������%�< H�[�~D���~��?��10�N"�hB�$�U
��T�_~UXC5�04Ay�t���"vT�q����V6XE 1�4C�ڽljMl�*��e�ѭ����c]�o�O"��u�#�&���/����ˌLX�S���������!�<�m�rj�O�`��M�],
��DSt��[��e���ͺ�����!w�TO�ɸ�#t�d*����Ye�k0`�U׿��e~�vཱི9�k/�;�e8L�;��K\.ȼNF��_�a�?WzW��	zH,�	^�u1Z%718������\�ʎFmÒ�XlxVHYEB    3d61     ed0z�� �Ι�����UAaPH�)�c!�1��l��g�0��ϹS��1�^$���>��S R9螜�B�	��$�b���a\�m��?�w\��s^�^GO��eX
� ��
�����a��$ɕ����Ĺ�8R���AR�D�޿1�E��-� �������RJ���YN�*�Nиt�G�F6)�^�gY�j>����oo�+	T3��(�I*��ۦ>�����Z�=�&T���N(��&R:'����h��X
�:��:��z���CĠ����њ�F^����D<R��E�������\\�;��{n�Ct��g�����P�["�J!�b������QDq�)c;�� �M�����	/Wq���c?Z���c?��� �<�;&�����W_l�{K[0���˽�����Ee΢pMAa���>�A'�)��\�WK�M��㢛���X�d6K�q���ZbFi�U��w3��~G�Qha�&0~$LֵL�$P�f�.�ip�'���1.zḘ����T`R��U9CM�3a���F#-�mxM0�����J�#ֆd{�tZu��e���@�S"R�EU8�<́��	�?A�`��G����Ѣ����˙3��~�1����/�^���b��8
��a�����Z�_�N�N�^ˣ����#�×����A���?����Θ�w�apP���[eY�� �yݠS����/�餰RZ��>�Eo�����(��8/�&'�K�@�c�0ͳ�C�O��"0��hm�j9O�:�gU��=ް����&zv��кyIx�3��_�"��Ėu}r{������i�F>�ļ������!�vg!�b��i�lU��YКR���y}��c�~�e�>�����g(�K����PE����n�g�Fy���ӝ�i`d$m,�֗���s��l2��ȴn��2�"�|E3*އ�,yE
y?�n��0�*��,��Ęc�I�� �N�W^��������&����e`��d[Tv������佖;���Cbe�-��]p��G�\����U,N�)j�������Č�u�R2�4�b�*���V�Z�'o�"w�u<	`;0��Gek?�~��+F��0��ɨ�$� <���ޞ>a�nѲBnuC�$+�~�mŵ:'Ic�P鋃��	3(�z5IB	�� #i��x�U���6�KF��VU�6R_�m�ct9�)�	hu��D,-͕��9(�[2��*k^���k�-��N5�$Ycp&�h���\O�,ǘ7#�#T�|N=]�'<�a���_���Iyz�*B��Tϒ��c�纟�)�5�{��)
�	��W�����K�k�M�fL�~ɬ�
f˽���)��<��@0"��wd�fi6�I>�(E(w�a�)��d�D���˕���0�k�l������|ש��I��}�ܽ=m���XS����p)}0�.b�C�²2X�} ؇P�lp��?Ubt�q8p��Ue�'�1"���%��J��
,;�
��0�u|��F�@ʪ���'N�%y�.�t�?Q8�ׅ�����@��3&�E眗�V|��'u#�Gn���������N��\�"-�!9)G�����\8�h���@��t,�����G_N��{�Mg��]�w�$����H�o�L�2K3�>����F��1���ţ@�?#O���=�sP�DE�%αj9m:L��Qg��{�|�[u��fw3���W�E�8)�d�f����+��w�&hC�]Y}��_�A6��b	:��?�c�N̍�(v~Pg��>�[��e"��%�h��w���_N��t_��pk�:��"��P�V�=Mȏ�!�R3?���2w�;��H�+Yʯ�r�`tun�^Zoa�Kw�]��K})��j�Tފ�-�w��͹�>���q��:	����0PI�3S�6	�Y�q��
��	)�P�+���L�.-��'�꧳������;9Z�=Y���fj���H?�LR�Ô�S<X�tWr�ĕ
�O0y����RdHۧU��Lx�3j��lX��w|��_4��>�u? LeK�g
gS.�v�;�������r{�����y��{�����\�,z�I��T��`/��5����,�V��c$��8���g����9����/�[�5��6��6���g,)��5�4�d�K�èﹼ�}6�HD����߂������(�)�>��#�A��hj*��y0�v��C(Z��+7b�(��K��Ѵ����M���7ht���
v�a��BJ� /�C��O]A�d�ޛ�"e4�����Ц���×��V����4��j�E=o\��m yZ�@6X��=
�l�R��_W�:l�4-�5��":T�-0�z�n+nƄ�����keCj�����kW���yl���.�D/�xъ�$�!��n��� Z.![�S���^�G9��y���B���&]*���,ȏъ��e	嬇�6(�;�/��E�%l����"!����{����y���B�T,g &�y�J����hl�Q�w�}�
���h3"Rb́E%oW��ڻ�HO�:Q����.������r&��%I84k p�$�'�V�+�&y�N�� ��%ؿʿ$�\S�vH2vi3�"|�CX��yc�D����y��6�]� �!�O$���Aoƶa�i�G��/��n4�3������!8}�܂EGH�n6��s|��Q	�Ƈ�l
l�P(^�Wꂄ�"�!$�yo��K�r�w�1/���6��0/W��J���"U0&�pw\]ֱ3�/��.9�Q���J�@
�E�zd�@VC�b�S�n�������VT�K��
��bR���w�Fg)��@��S�X�f�M��K
e�����5���[��sC1w��zj��$ڣ����)�#wu�6���_���G�)}�� gK�}�O��o�Z�]�κ������H�=���g��������bD
�Ҡ��e��6�~0������t�=����]ؿ�*�o����w�-��Ŷ���9'	u�c�ڢ4�h��A�>{vji��8
N�b�`�2���-���!�8�(/�8X78�șm'�0�˭d0�q��jc@MK������dQm��L���5�����^iK����;���Y�4)��9!3e�Ƌ��Ԁ�6o���p׏S9h�NV���r��g��j�
���28�VeeǴiZ&4�lLAX�DL�������&An��yJ;��/I��P(2X,���.+2�q�O�����r��Cz�' S�O��P�����`�7T�kΕ���#�p�O����%�uq����A&r8���!�j���>l�����n^�[�<"���:��Ŏ@����:N�����;}�c_��c߲F���sˉ��6�h�^hqgS׍�Ʋ4�{wvBb������� �� ���{$cJ5㮁;�]�5��7�p�]Vx��o��M��6��Ê�8G�~�`]��&�`�Ȓ�<�򄄏́�q��x�}��,(7�Q=j(����ٓ�Y�"9P�f@YH̦��z�6u"[�1_�h�U�Y����d�Z�D@(+��CF�]�[�`���U�jH,��Y���G���L�˪T���54�<���?}۔�����!��X��K�ʦ�E���K��83�ՊG6fs�Q��?6�d�8
�����MK��nG��2��hy!W�^��̂L������$�)���� �K"�f;-�!�a.