XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���|j}�]`zZ�ˇ;|Q,	P^�X�'GO��i���m�v���d�F�4�jfA��H���}�9�f���/�S��D���nB�NS-F�v�d�����	GmJ6�������j�A���h��Z���4yt\	�ɦ��;�o�"��%��9���i��E��AP�G6_٤�K�VVih��Ð[�9�T��uP�!�d��t�����Sk��>��� T|H�x���Iq���C�#�mѧj��A�-;$q�����\
'��
�A"�9�9���;9kn�aNjl/��`���s��5P��c)��ZO��[�L�/���5���d���u��� ��1�B@��&+�ډ�Z�@��|UD�Q<�C�{H;̓�O�(����Ә�@���`���gK&�"X�P-Y&��������y����0"�w�x܀��o�9�TG�Y�� y��ω�K��+"'߅�?0�̀f�p�Q�ġ&�ь��G[�@ұ�r0�J��Ij���x�\��=_�τX�I���=�{����~�?��bW���c�H�`d}M�M�'M�A���T���#)�	
#(�4f�,s�r��I%w�@ե=Md�ѽ���eGKƱ�D��}v�ΞO?�}�$2#?ݿ̮$,7�R$�ɳ��|4�,I��H���B�V�Pq��Jh����Vg�aڷ��	�ycge��� �qԀ �I�ő1�����),KɵBc����'ZKNN���a�y�����(mz$����ܰVj�������T��XlxVHYEB    fa00    1950i��\K����ʂ���:�hI��J,����*��vq�y���y�\${��s�W%Ԥנ���p���6h|C;_��{�!������RO�?���|H��k9����5lJ�����:�14�����>�Q�"ZU�s��r���_�~��
�N��m���y��pl�.���J�t�E���&Te��$8�u���v��[G�����~�;�O �¨���[�t>���J�}���Ym�A�t0��c�^�c�%n$4-]�l��b��q(F}Qp.<Eq�r�>wyy�{��3�vL�V�Qk |�J�X�؜�c\�>�R8�U`O����2S����+�[ �>
���aM�������Y'^C>�x(z` {K����'l�Q¤��jK����n���"4���qϚ��}��s7S��Sb���ث�<�y����:׳6C�"| ����$������l�m1N'+8+�)��8�w5���Uî��)�Ȥs���e��Ty�9�(�|b�H&D�u,� |�5O�w@�(?|�?�i��D}��F�O{�
�����[Q�e#q��p����3�-a�*r�6�Ü�"�Tr���n�s��/.��;Hx+�Sk6�md��?|S�TJ�h t��E�r��:FP-M������_!'h�[eA��g��}�����-C�K��c�����#�饯W3'�S��ϓT�p]��wԵ�6��((����Dmw�EzBě1R��T�i(���Iď�f6��;�!�(�ۜ�G�8��P���T�H����M���Շ)��k�k��;�8f��:���Q(�� r}�<����e�/o���@�1`����B+X�a�L�29�2������wZg���&�ޟ�;���>dke�O��I��3�������8�N%��h�@��9O��I��nN�w����*���d��݄�ʹ¼bo=���g� ��Þ��H�*��􃋨�@[�����`���2��c*����m�FQ�Cs��j�Pvf.w5�iq�
1$��&�W?�0E�^Y8=Q�2��r�a>$A�G��u2���a:Ѕ�O����	-i·��| ����ц����Yx��N��h��)o�����P�Vf�e}�r�����)���N5�9�l�0�� Ũl,kY:�ʅ��66�a!;v�&:���URM�P^0��������̵Q�.��P���b�qð	qKICO��$Y���&��IL�Z1*�U�qYo��+�K�w��Ko�f���
^��
_�T�k][O��=��઼_Ћ���0��Ս�|4�!���<�oyv����(Ha"��F��teuz�=ufJ����W#��_q��N��o�0���K�)���R����(�R�W�_BG��H5υ(�S��.=�.��1cw��>v���Ǉ�`��ae��~y/�WI&�{�g�0"�j_<Z��D.��\�_K�i�8��߽��C������g,���y������/��0W[�@�CSr�"[�J�Cgא:�����B�g�K9����!Ӏ�ඎ������i�H��̸��ި���s����`rs��c�؉c����m�z� fsĭ]Ӯ�7l�H�,_�F�R�i�h� �y��`%L�0��՘]��P����0ؗ�I�Y�ovٿ��;}���j����Q=��a�ey�F����S���, �jf�k�8�bK
p^m	���o(DR�p�l��T�<}�|I�B�*b�8�KO� x���ږ��6�7�^ /
�%���3띛,��.��P�����$�����5us�3D6e�z�*�,��n��irk)�GH"�Z:e��ޝ�w��X���Fۉ�l#�'h��<���_�w��T���ݕ�=��/Y6B�Ԑ��&�{��h!���`5ˆ_��(�ݏQL��#	�w d��X�xdÂ��(p*uY���j����� ��)��L���"߮J��AE��{�"Þ�]�v�Cu�'{_������k�d�����=����d ��֒�c_�+l���@���O:�D`����[��}�]u�Iw��K�H�A��*r�P*���΂m��!�n��G��W�����x;�γ��!;�?�e���h0JVߋ_z�ٹ� �U��;躌h�V�4��A��wЕ65Dʔ)us�"Ǯ��a�����V��=��@��,�C;������D��*����#��$)$��S�wf!�z9�����j7hy��� ���LVS�TMp�Y������@H��lUH��H!����7�M���#��H|���_�2bݾY;��r���`�_��oQ�7ǥ!e�dna�r�(7����y ��a�i�y(�����+�M�!�<!U�u�sZ�'�Mw#2�H�_@�2�萱q� gy�zI)V���h�������H���*�Z�m�ݖ�$ˠOl7�y��:�8��P��@ɆO&�zf�)�*�ۄ؀�*cS��Ym1��O6�Y���/�^1CT#P"c��E��S��b���(0[�
��)3��Y�e�� _�����Ԇ��<��|���y�����_j���jo~-%��_Ň���r�r�;EY#|�d�!s@��%Z��-еe�m9�ۨ^dZ��B�|�&�4�$Ǳ�6j��Ggr��C��Y�I��eDK���8#ߟ��8w����w{;��.�o�.A.jh���/�)�Z�	�+���)�:�g�,��:�d�-ګ�	����S���Q"!����A�����CD���J��Okii�rǔERkm�!���u�3�`�k�}�T��������7�1h�+U#�j3����;S*2�:��.�GI��AAZO<d�/z��f�sn��&�KǾ3�δYNġ'8��BjjX�UC�y;�n��i���#���M���K���Π�n�{Z,`41��OO���n����\O�@�����Ea��2S(�u�~�ɿ�s��o�<�Wzئ$��_��M��&���	.J��T\�ҩ����1�|Spp�ztV�B���$�N�h(=B�l/�� ]Z4��p-��:Ƅi5�Yߓ�r���y���
B�l=9&�Ro�Y��
/)�OPͿK���M,S�E�p��6��HK| ��2�}ʞ�[�XG:�� ��ɔ����"
�N� ���_�WHщwo��?�XN�8;:�{	�ؙs��%FF0:�<5rʻYDB�٪�~�n��o����W�<��ǒaX��i��`V��j��}��䯚np�U�T��7�#���r��&��o����w����[�=ksv�8��{4[�2���L��S�'c̚a#�����M�İ���������'���!p�)�v(BwJ �m�p@z'��(@;u�J�B
+��x@��� ��}�b��M+b��ۊ�_��D�d�m@YꀘY�L����v�ͺ�cRf�2��_N{z���jZx<����)�����šϳ��xGBs[�ÁuY�f�9P %�;�˪6���-�����*9�]:p��5{g�8��ID��5>54p�F� U� R�ص�Kil[���1���}W�P��,,F���o�h48M"���
Xܥo}�򠒋I�E�o��\������}�h�Z���M���B���	O�ia���ٔy��={�^���A���[�J��muB:�z_C��^w�%���,l2��M�%����������|1��_�e��Xg_Y���;������:��jq��)K���-x�Jk#E�h��"���G��`*��9k����i�Y���9)�v�gaL*���	7�b0���h�5���B��[Q�����8�u����~�p*5�|Hz@یĩ$:@[���<�ǒ�N�l9�������;B��EUR��IG�q�$u�����C�gH�i���y��6���g'�!���irGN�*�"�Ʃ%u$��k�T9�1�A�ƞ�(��u��(W��.�ByE&t\�~BP�bnL��&�8å�9�R�%��#����������i1FK	Pl����I��f~�zZ)�7Cp��T�E�N��p� �����/��8���f ��7ª��&�0�$�a'A=(í���������3.{r:�:�q@%	 i�8�/�����T�]xA�ɰ�:-�)���;��:�ײ����Pr}�l�c{c��x�V�ՒW�f��+�}��4���d�>m:#��bZ2��!�dW���S�DIƔ�i�'T�̓��(O�}aDL�btK�[��O�b6�.?�C2���q"oL�o���ͯԼ_��Vg��376hC�w����
f��B@\�='G��_���Tbg��`1t|
�3��pŢ�WPt.x�)#A���`9&�J����V�#�պ���W�l�+x�!J���A$�C�P�1�����G����:��P��� .������s���%���W�`sٮ�����{���j=���ԨS�t�f�I�r'+Y��C^�b�3*�U�m�(�g�m�P���U��
vCݗߑޗ���WVelF��n� MCM:�X�8���E|#z�����3sdU��i���ޕއ�<q�|�� �=ɉ��'x$;Y}�`�=Pʩ� ��=��s��.I61�_\<�� W˫��Zg��Y֪�5�oWs|xqW�
߸��F��;��U��d]�7�>h���{����mc_��%J-��v���b�1Ϯ��.0�۰�+V�?N\�d�y���ğ>�SZ��|�\��N���o���: ����XjE�R֢���\�N)��X���j(��.�`��J�@��G���
tI���t�� ����^��,*A���b�).%V�H&U�����d�q¾H1��B�\$��͚��Y�$�[�[p����4�.��`.��,]'�����܀��L��t�
�m��v��-a·�$^Q�\s�LKf+O�yUd��a��G�y7Z�+�W�F�A�@Z�«����ݛau�hQ��|�kp�"eU�h���Ӗ�9@�A�᷋��?���pko�d�������+HPG�Ƿri�$*��+�Zn��4�m|'�0�b���|ʁ��	EޅSe��s������~��06Z��Q�v�n���:�AF8��đp�����j�u�Y爣ɂ.d��2�"�"֠6����#!bx���#�/���(�����0�/(��^�/9�������]�~Q�����^ �.��*@%�h/��K`>�W��BY}���~��/�~�h�U�~.�g}�ɞ�e�Ŏ�����dd�otw��}8��z6�.��z,�����!���ȳO�2�X������3���Y,�������'��U~B3��s��>��*���*w���"Ar&�]>޻��X/��q'��G�D�x.�"�4�xIV	�6��B����D;�:/Z^�*� @��l'�FU�+�І�6�6��5�7�/�� ��J]hv�f�7X��|YO�`l5���]V����XL
����= sx�V`옇;�� ��d�y���=V�4�D�y���1�<��0��UM'�`�V���7]!�vs^@����a�s�ur�9"�԰Ńǯu����W��Z�����)J �7�H�ҍ���,����������-C1©k`+��5)�ĳ�!7�m��N>���wb�b�~^��~�E��X����љ@���N���x2M��i��r�#�Mndd#���ɦu�
�{��ȍ�u���w6,���m���:��I���X��;��3c=���B2�Ei���$�����@��ҙ�#�$����ٷ����I�L�ƣ��`t�Qݲt9����pJ���9K���Ԟ�}3���R�n���%<�c׹�aZ���GIR�9J��!H�[��;��tixN�q�;ye8ϔG�U(׾��H���0g+�U��� ������t�q--oV����v�<'�9`0���2۷J��v;�g!f2��h�a��/[n�0D��c�Ť�r'@�X*݇Y�R��".�d���Ɨ�ۅ~TN��ÉD�o�	Z;(�S̪���������&x��k�ǆ�� KV�����;�� �e)u}C=����i̙�d�V�\s�_?�����F�}x��5r���q�?������ꖡ�{*�1r�0qi��$C��1���'�g>��X�M���t��#%,�g�5�2�!N�
���q3����-�`;+�%
-Hu���;C�=V�jW:�?�F.�w4??h:���7��9l�hw���ٔ�K����{�������ʬǡ��E�*�u�I��/y&��j��щ�����;��œ��!ӄԚ"�b=�3�����Z�^XlxVHYEB    fa00     700X��b$��K�	3�iL����e��1G��A���څ���41�;�Q�mI�Q�\-9<S;Rg�H�UJ�	%�y���8�&�O�N!7�]D	�Rk��p�2 {;e��]ܖ��Yac�+N6,X;n���2���*&������������)|&�nГt*4�h$ƚ�;��=�;�=qr2� �ꓩ��!{�`b��X�Y�~us���w�\:�r;+�tm�S��-B�D^UL���v��,E
9u3y������#(�K-�Fz��CQW��y�F�9�`&�&���ޜ��04�ǁ��7�>�퀙rS�aOc�`)-���=�P9V��{e�4)%Hi�U�Gu�$��@3��8;!L�ʛL�4��)w��,°� ��T�5�{d���֙��s���2�ݩ\	��{�]� �U]���r�R嵉/��&�u5ʲ�4Y�S=7j���ɟ��@�Z;�#QAb����Z��Ỏu�l�&{�s�!�A�d�<��"ڨ������8����P�D�jj�Pp���.?4'����*�9q���L#�����b��W�O��B`kv�L�N�ʂ*i�v�ʙy���a�[�W���Uz��L��;���#�H��5Qy�|8�V����v]��0���Y~�9$�o;�<��S�`� Fh��
�W-xFN�5w�����r�V�@o����.;F�v����Q;���@��iF2�(�E�VUJ�F,p�㓎���Ge+��_2q�����/V2�.�^�I��_G�����`x����FS"����ל�*UcU�.B�o�Ą��ZӵC�r(�Ɏ����X��O|���Z%!��3�J�����CFG��و��M5�6D���]�ɴ�H�(���I5��)
������ݸ9.p���t�A��YL��Q���)��F���t8�#�ݛJ����I�MQXt�_h�ؓ`�jL�J�� 	�*Mw��mMȰ-����_
��n �?�������p�������EV�HȚ�7�.$ʾ��}za�q%�,Rr	�RmY`ZS��b���R�mb�0���d6W��ma��� �
98��"�Lb��:_}Uy�u
��K���"ʓ��}�˙�:f�����U�D�ϸ�i��C�	��j���`Ȧb6��$٘���8�K�B,؄wLǨ�G
#)�1 (���bf�j� ��-�����KU��i��`��Phg7�RrN�*�;��Lh!~�L1tZ�X+G�)�8*����)S��Qj�o iW�R�Ĕ�𻷛�0*��kMPV�AwJ�D~ �z�����bUt4�׏����X#�5
rkO^�%�[�ȅ]�8�i,���/���/+HƁX/�?{�,<�F��8�*K�3w��f�b���ƚ���s���^S��x|�]�I��3�Fr_e3!!DH�*�fsY.=t[�kDM��N��8���.�i���a��$i���S�
��*��!�\_ !��e�u"��
��^��*��t�W�:���x��h0b���X�/j���c¦��2]/����`or'�_%`��r���&jy�)B��2�!�x�E���{�-���
_��Vn貽f�5`X������"d�T�PXW+Z���)x��ct��7�Ѫ����kc�P��aIs�ח5z���`h,Պ�W�6�M�`��oY�]��{5~KT�+-j�b%��y�9JSD���|V�� .9/�$�"�{�M�7�-�ZW��K�rk��b�'��!0��,�������<k"�?XlxVHYEB    77da     a60�-S���J{���9(<��Zw ��m�Y��)���.�틨�����W7�fd����&�3���Q�ƙ�J^\�5Mz�+[����A��7�K��mA�Ӆ�M��϶�K������$�8���jӁۏ�,�U	N}����=���ݲj-�:��ܶ+�\�W�;&�Ȉ�OY���Cq��9c�}��m7Q���i;�#���lG�I�;��홇_o��#d�����O�O�����w	���5eH5�kXW�>q�i�95���.ZpN���0��I��A<a�Z�5���T�`i��Z�$�ej����_���O^���ݛ��E	2)���U�>�0*���SIa���P����]���w�5Ev~�r+Nڰ�T���%l��9�
�E��?�y@������j��͖�C��+"5�e��G<�����YX��˺��i�e+PjHpS��L��u���MQ��N����A���}�
��.�d����;�ک#5�ڬw �\��O�_H�:ĵ��7j=՞ 5�S|8G�hk�E�g�a���b�b��g9[�x1in����������'����q��rI���; ���]����}�����EF(zW��-Ea~a�}��R!���5�I	w��n_�x��T�1�P��fI a,^����i^iq;�/����2��CD�D=���
2~%U�wc����%Y�
�aF��
R�i?f1���f�$2&���Ж����)f�Ѧo-m�O��u�2��6�Xz�] odu\B�pg9�J+=��u�s���N�&�Y���M%S�Xӆ�fb�� _`�e�U����D��.��Ð�~���,�s�FP�������#���5J���W�f���5y{ ��Th�9�l)��?����&�����IJ��M�����w�ɻ�J j�;��N!c��𲪙$TA���~�� ���*L����o�_(��XN{{�6wԁsj����ؤ��f�����4�۞4�z.�H\�
�ث���%�(R��1.zQ��HN��(�}�\�M82I���6֨��V-�P6�}���X	Ȱ9��X�p�h"�!g����Ѐ�[ mh ��瞊��C��6^�Ǌ�l�V�zWt���KXB�lg���r��F�X��7��x��k�Tz� �n��u���S�5*-�r����~��dm#��%����@^�9>�A�?��c�E�NMQ�o��\�B~��P3O(��J����6X+�Z�H����6!��m^W�!���Kf�si Vi{˻�G�RZw��=9���Up��1��I6�2A�;B-����x���R�bG�t2���;�*��:� �d�F�^�u�3:�%��<_�ߢ�\�|>!�'���|t�ש�����t�0h�5*;N�<���SVZ�V�� vĄ����c�ʢΎ?F-w�=5�@lW�;Q�[=��V����ڰ�(H� ���-�����FX'�i�Jb��1�%%.`�i��Oq"�"6������W��
yz�����z4�����HF�~Հ ?�l���o:N88�9�I�\Nnx�}�3#�z�

[��%��f`;K���˘���R���s�w�ͫx�	�w~v�Is�8���� ���|*�7��R\�k�B�R}�|PX��d)5��Ik���&�/'^ �"���H:D�P؃��A_�����]�k-��+n_ذ����n�������]�g�d🺄�F2�������l#<:�GQ���+}�3K�XLj�~A�q��52+�E�����^�2�G�g$sQ���ܳ�d��X� �]o�P��
%7G������~�,�9�37M�%���[Է���P/�`=��gsf4��U4���Ѧކj|�׮�A��A^�������4�C鶛���$�4�cg4���$Z����E��Q�	��k�S>����r�j�˖ R&nD�;�OL%�+w(��@��(���'F
��o25ta���y�!s�I�k33oD:G�_��6��WV�ΠC���:�rm�ڊ�8�t��1��6��E|Ȇ�?&�$?F��o���S�'�~x��Q	���2�b�бr. �������;W"�W���fA�O]j0�������l��>�����RX�ܓ�~aU�(��K�P�3wfCP�k7ÿ�Ɋ5�<]��:*̌�>��U�և� ��|�'����$��&�G��Z�h����%�+���1�	F����;�5Ho(��$B�U��ܰ�,����7@K���\��Xʴ���L�L�G[|r��0�h3�A��_.4�����<`��-]N�mH�����.�I#�ޑd��;\��|�O��H.��Y�� ���H�Z�S{�Y.q�D��>'H��ܔwϥ��;�+�1q?��qF҉��IV3��\B���[��`v��{B��A�t���x����N�n�G��7����I-N`�^j`��W7�^~qehY� ����Y�}C2��sl3^T����=��{�H��蕹[.�yűk��߄K��&�T���%m�;QS�t�����ʛQ�K?ǧ�aSVҺ,q`�<O�B�w�����р�Rp�F�LsF