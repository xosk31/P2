XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��~��57h7�f�;U�Hh C,�徹�{�b����[nr��h�b �
��6��}��>s�9��^,��X��U�;}�(���<F����b��SNM���ʩ���ec��+$����}������T?_�y�K��� 4Q��k���d�ac��I��o�ʹ2�4��{�wf�����A8���2@
��Ԝ1!�.�f�.x[.�+����}�fț��0i���E�q�8ѡ���-{�Z@g��B�<�Ľ��Mt{^}�OE/ކmJ#,�)�wZ�ͤ���O� d�D�}�N��7]�/4� �'a��(rz�� ��.燚���L�}�7`��2�}@��"�����#�U�fT���E�Qf��}/��P��C��[$����ھ�@� A��lXc���)��b͐�3�籪�����@��
cc �/��C�D�;tͯe�6���x^��*ڣ6��P�P:�3����n������y��8.9��s�C$�!�����E[nu��Q�m�����w޲�C����DM�q�Ԗ����'o>AD�c����� N�3���DCO#���Q��4��SA���AP��ߌ�#�r��u�5yہ␪�������@����"������3��Z��pa���c�5�~׀Gb��*�����~���N�f9'�b��(�D�zq+�縩�����V1Tw�P�.FN@�9
:�����r�%M+����W�Zv���14o#�m��~����(������h�xXlxVHYEB    6cf0    1960�&Mù���
�]2���_2�� �����n/�0�1q�fF5�P"-�E�i�7�~�e��d2�QY���N�@�`�/.��+���Ο�����yN4��Q�C��q�(���� C�{h�����VU���k�x��H��^�b��p�s�����}���a��[�������p�4�rnZ�s<��!�k %^� f[2�jzD9�`��!��WU
�؜���� Y�
�Q�Nd�C�# ~
��Am_�1Q��e?Ĵ{��U���`J�Uw��.POO���x}	���#��b���9w#x܋���y�H{ئ}N6d'�!nz�)�ߐ�;���z������D�RJ4�)��~}�8gE��9=>Jy;��%��O���&@RuS�jj0��9o}�ށ�`٤�Vh��+a����8pL��V����$3)H%Î,��]j�}!F�I�����-`��d��)�ә���U��9�ʔ���� �	��6K��q{�U���+P�N�1n���t�}ߛDI�
~L������j���$��lFcPJ���@T*lݬ��1n�E��%�X��Y��j��M�y�#����4�R+�ʓO�{���=Ƞ��r��X�@���g\y��wxU�^���p�	_0���Y24�)ҹZ(z��r�~OM�A�Z1��B�r碧H�^�Sq��	������=րx���;�������_�����Ǔ�)����2�p�:�k�v���[$��U�Tj���鵄�A�5�!-��?���T���\T�sԡ��>;O�� � ���~cl< $cHf�t�gw;:n.F�$D�%��c~�)�"H+q��OC�Ma	�Q>2%�m��Y�"RyԱ���軣+�Vh�-����i��gn�"�����U�\*<��R�wG��s���Z����Uo֢U���i/AX�L���I*'1v��G�&��EgϨ��������KEGx�����QX�똊'�.mf�-���)M�>BE�\�h�~ߣEaFCm
x�5 �<�>����~�p`_����r�W�,�Ьƨ����C�Hx�rfm^�oW!�[����N�['S<�YA���x7ca�j���OU��L� Q�o�Δ�R�� ��c�p����#L������P$&gq?��]fR����)
���5Sh��b�y�!:�U���Pc��֓`V4!�+�U��M[�1��hrZ�p)h��T�~h�Ru^�*��E*��5\���R5�D��A���?r�;R6`����Ê[�0��O��G�+�fݭ��ڷ�M�7칙#�h�_ �F���H<�<��8;X�1��i0Z<��j���R�Ъd�����L�9P�4kC�֩���}���A֔����K�"��0r�=�n:�t.��C��P�V�ƌA]"+T#F��Aj�w0ŬL��^�&bZ���g򕴵z��r������dZ���p�lZ/7�h��U|�*f~1���+n]� $6{6�x��.�ѯ�3�$ɒNvX�Aci���v��X��d爪��o])]�I{.�N ���i��@[;���4��W��A`�"�L��Q��wP}��d�k�-\|@��;B�C'(�dos)�d� `ͥ�~*N���+:0��ɚ�����ih��Ł�����1�����F�l��n7�$8Sk��J�����@X�B���PU6���\��DA�)�?�އ�P��1ot2`�u�V�tDf��1h�،���M��=�02E��*�ߏ�j����P���z��J�V`s�	��r_����T�^CW�����%�V��$��p8`sR�nX�I��z,�q�u�~����JVh�+���Ӫ������Р藘�(1�a��t��
���Gǚp	<�$Ɏ���,P	Ž_O��f'��,����d\�8��DO�rP�8h왘>J�Qv��`�����ϴ�����'�v
1�(��>��&���{����׈���rlr����� �wm���o��xת�Ы��k�{���[H� �Y�3X}����f�i�Qt��.�:]3���Y`��P~]� �εU�Ǔ������]��	^h,��R��.���c�����ª�Ȫ��C�4��@�0�Z\p�qF���wd��c��րo����I�-�+�ln�!�f�J���~�L��-�'��V���X�E\$���^���@��Qţ C�-���`)g䂿�Ə��+l��չ�ԪĒ�ΟI�hG4\|�CB���Ƅ	�w�پ��f~ƹ�? e�b��)��~Ood�K���<� e���Cӆ�$�P��˩,5�7�N�a1���W�/��a-h�${�����_5�����)��Q�J��,z������B��@��Pt�����&�PoXBH�n��s�t���M-s��������ڂQ0�-�w{��ԓ_s�t��1�(_�O`=O>��VZ��^�1����c�lT�0�����t���U ��A)ZE�W����m����2D��<-�C���x�ee�����Z�R���>���+���J��^���E�O���޷��:4����߯����o�N�F:(�̏�H�Z��d#�ݥ���y�<�����	U�[`�j�ȪW�x��:fa�0@�@�m�[Vt@X�����"A�Z�&�O"�eWP끛@��ި�ry�3.�y��{2�*���N��)\�y[��V��)l/��
X�NfuB���A�8l���m��D��P��b�����V<� �c�����YX����h5g�;��Fڋ;���-?RC(ģTO;o�S�ϔ���tK�ʖ�-c[0�F~e	D��j:���F/��E��D�~h������ZǀSj��+ƅ�cȯ=��bE(��@g�`����UA(�9�z@�b5�K��鬻�2�0{�[�?8�A��ҹ$�D���U��C����'��bK���,s>#jn�`7Sp�2�f�6���ҍ��{�Uu�$Q�	����u��� ��dGY� 8تE	��G�i8����g��"}(:���b'pc��������{��2��0���`jL����kC���q���;F�'����l��z�����G -b�S�~�ǒ���9���7�(�oM�A���$
#X��}���)��&�'JB�~��5���Z]zkz�[O3����m�r	���B1H" H�v�;?=d�IX@JK�,��"3Յ|q�k�-e�bp���^�q��(�K0���h7<���ie�ٮ�h�麔u!;nջ+v�9'�����Ӹ1�0�R��������AK��>MY�9K�kn]ӹaeǫ<��gDQ���h����x���މHf���D�5�*�e�u˙��^�'~gN9�"��_*2�B��:lΫЗ����Ŏ��X�/��s*��O����v��@х�^�FX�4v��=�<�M1Z�ٛ�R!��R�����f�k%�HE�Ӊ�@ϫj2��/?�S�5��iَ�9���K��e�������0�֤�3���g������ ��xM�A�^|�
ʗ��泅?���}�Q�F�:j��HK���+�U�q�{<�D#�Qy!�n��os�]}{ �Rh�k/���	�ˆO�R=Mf3k�w��|Ml�� ,%���zl���FM�8�ygA�x�p��2͍��n��^|#�g@����T���wf`�=6�3�D��wo��c.�4���{�맜���kX�c�����	���f�`/#���むZ���T5=!�a��8��ːi�q�M�Y�M�V�w|����
���v7�fF �J���hb� 9�Ĝ��O�S����7!������@?�+pǋ9W�
[�*�U�fg��~��� ��&�z�Z��΁��T���0��[��=>� ��0�y�\�ĤE���#c`������a�Y1<u~'"���#�:�� p�b�2;a����;G8O�j4�����A�����]
=�p����=�����,G��E�[WC}d3�R�<�.͌��ȭ��|o'Y]�h��X���օ��g�_X��Qk��?IY��%ħM���2�h�w���7����PS��X,�N	}��To	����˭��J8A���87���`3$$�L��Jӓ�XqM���I�U9Y�u��ȶ���~�(�cE���1D�75 ��MC���k<Lԟ�b�v*ÿ!p�N�-��RCDsL���*��T-Pխ%������J:�i�sZ%8����d�F�ڈ�m*I�uF�܇'OE�S1�	.,���Sd�s�Ch�Ycº[�G��@��u>jf��mN|aܰ(V*t���dv����F����`x߱NB��ם��7�O,�>:h|��l�p�����~�RGNP"
yP�E��RɕB�?�S`~����2b�wf�ĲK��Q�걪i`��`d4%ϗcɠ��� /Y8�,�M����dS�1��ިO�	�<�]D}��q��I��q8=���`L�{,��6_�q_��ۨ�%�/5G��<q$�a�`����Ҵy�N܊�� �+�5�}�\�����z\h�'�v�FF���{����;I���q���������)M��	U��cj,(NY�r����X�P͔�"��Bi�
��PnҤ�C�YjD���Kʢ�(���jU�x�/���bf�i����8���r��"�/��-�*�s��b�kus���^�!�=�\co�-�W��KM��Ԛ�QYo���k��[����n�
�!� �����Q)�_FW�c�������5�;)0i�j�!����h@D_چ�:X��7RrV�_�P-I��L��e�0���2�hcL9@:���e��-YnW?������iT$n�Y�
SњV���n��m�ţFM��S|'�/s���ɻ'$���L�d��7��<��]�*2����Y���`2�E�`����Nq�֣��k�,�3�/(.����46�wO(�@|�ɶ�x�Q�)=:nm��!�4�����L�9�"4j6|�i��P�3��L���S�c���95���xP��'3{Ԯ�������ǯ,�L��*'��˺�q=�Ų�N+����]~���P���_!��k�l�w��Bș\i�P�����`7��9ˊ �v�;���VM�xK�A�EF����EB��c��C��j�?��	yn�clO{�w8�C��$�����=�#���{$��"��l�#���q�r+�1����Ȁ'9@gR���oL�;l�t���b��CzȦ��J��{�ءvCOA{5�a��oE����X��~��ՌN��+��%a�n59�l�N��G�����
`��X)Q�bA��	L[��ڙf�=��E�"Qt��t�uEaf����*]7�Ib���o]� �h	����sj��	́�I��~�u�m6pC�7��Eђ�myw�JL"�j�b�8�O��*${J�8dQb }��)�w��1�����M��+��C$k���qX_K$��8	��KZ�UԖ_�n�C?�bZ�֓��"���sB0 (}���6�O<�k��n�C~c�;�h��h�t]A���V��xM�j�#��.۝��]Q�?0�8f\��>G5T;Eڋ4=My�瓤�f�����&��*�C�4��Lb*'�3�t~�~�6�v{��lM�O����H"��	����]����}(��%]C8;iW'��7�)8W���7�I���G��$foA@�����@�6�q���S6����r�'�`7(����Z[]�n\�*��q��E���`��ӏ�m	
o� ��)j��p��L�H��v�l�b{�\�3�_x"t)�3��hL�ȫ3���2�5��z�9�-���$�o�t�8]9���Dj?(�v!B���ë��M6�+.S����	��L��<8�/�{�c�u���+w���
�0�� j��K��)9�n�]�hXZ��b!I����{�'��8�z�,xQg9 X KHG���?��4u������D�{B��v��i}�.&O���A ��t��c�rvh�zHU/xJ����"o*���"*Q�Vn��������=���?�7�����2Zd�����Q��!��)v���'nE:.�wqfF�ї��^�`���:���"l|"���B8$'x�A�65�]��iy�g
)�I�Hp�".�y��FO�[��܇?��A'�I(������lc#^NZ�d=�
��<���*L����&RL��9V�)ԅd���mFtL�a$�Lla�]�NA��=`m�R��9\o{T�f.O��̓a����ǈ���G�l�=U����s�c�*^>�k+#���� ٢������о���PL���ES��wX'J!�	[�^K��bY�#.��6i埴f�jZ9�|*��m��>!�օ�)