XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���N�6c��@���|�0��L�$A�ܠE�5e=���Z���~������S���Uo<����En�ą@����X�l�R(�h~��5Ŷ��6P�qڊdg1I��(��Xk��O�$�%#�}��g��k���s8�I��J��&Q49�Q�ѪD�8��n��H6n�o0:{����i�x�_ �Օm��G;&��.| �n���%����ۙۦ#8}�9�Z�.��k�զsG�CI >�)�y��n[H�z�ϑs�MM6�H5�'��/�?7cjg]�\�_ʠ��)i���$\�%}H8@σ�K1���Y*��5`�'����
�s���p}���3�v���6�U�T��q����}Y�102	uKNǛ{o������IӀ^��DϬ"l��%>(QI쯻p�lU����3gO[��P�尧R�*lp}eŝ�4o�az2���"Ů��FuB��t�lf��`�\��5*N?���/��L�,��P[��JQ*K'/�U]E�7�j����B|�	C��u������ٴ뉬my1ۙ� X�O���;-��Pj�&N9���k�o���N"��*7����PZ!�^�'��^��������s���p��*����|%�)�-��j�[Ў�Q6�D��|f����+�34�
���P��!O]uT��i���?�������\�pT���m�֓2�D������$�Ӛc`O�;b@���RP�C���帲.^E�8����F0'R���KyJ��G�f6XlxVHYEB    2a94     c70Gcs�p����٤,��ͤ"b`Ќ�!1!"��S�I���- o������D����CN�H��R����D�XS�j�^�h�c�M���ش�m�y��_��0�_
�Ϡ��,�VNN,�0ޏ>ؒ6��G���?yQ��$I�ࠊ�v齣�?��J3,o�QC�Q �����u_J휇�!�o��P��ֹ	��󰁺�5{�KU��e�u^DQ�US��;�����w�#5���D�{�䴫F���(��>S��w��T�a�f�)1�����H\�`�4��A�����M�E��kL�M�䇘 �D/LRy��
>ѺN(�����LK'���K�b&e�x2�-�����I�����[^a�֦�R����̧����Z�}r��d����x_�C(d�^�.�_��;ɣ9T1��d�bȮ��R��b OS�-������x��F�˱��Bq6�%��풄GZ��u����F�M����0�8�գ�?Y�y��z �yj�O1����;���@����ۜK�dé��qm���ѮG��YU{�^WL����p��������$�e%0�z��c��Q+����=.w������\zŵ�1�U#�hb����;��F�F`�2���H~:��2�)JBT�lm�/�����p�S��V��\�t<x�TrE=��y>7�w��c	���zz�<^����j�!�'f�;W+7�����St\	�)�Y�n�ĝ�خ4���4���Z�����v��r/U���:jܥh��ޔO�N
�hƀ���Jy�ȣkU�c^��gt��+~;����Z�����f��Q�t� ����߱B\�A��a�v�TCf�������n	�x	M���&|�z��8)7�{܅%{��եdq�Pk��Q��M��,���
e��r��uԉ��C�����J�<�a�����C�'J/d3�6)�Od蒫����c���Y�����S�mh��2�JMuRY�s �M�?4�H2�7<�CpR�[Z-�'��r�������e/�Q���aJ����	\�G3����P��O��9dUR���z[�L֐'ƹh��vԑ�O�C�f
+=C��SHc|�S�V�`����v�t��l ��ɯ&��
쬬���?Od8���l4hj�R�m@��o�i���V`��j�f��u�$��͚4z��l>kў�����7�H�M=ë�dљ�4e�M�#C���VUjl4��|����\8^�R�[%�H�"���M70�*�j90���f���/n�WꍾF�L`Vg0ga+��,lY��q�UTD^����\���]�"*������x)Q#�ǳ�`,��S�vV���R]�8�6���ΈW�!URCŇ]�n��r��%��z�	�V��ǧt��%J����=��ƅ�}(��V��A� �����&Uzx���av�Z���I'�`)q��:�!T����G9���k�5�9�<]p�~����'��R �(���	9g/�6q�)�H�|���,oH!4ro��\(R�}|E�� ��H��Y�S�@h�A�&	gE3ݰ=�{<�N�ts  �@A�8�Ҭ�M՜��"�.�,Gㄪ�y�uN�oDA.�s&�k������lH�]}u���J٧�@i$gQ:_cXj���KҰEǊ��[�8�ބ�X�b�PSO׬�~������ɧYgC:�,��X��<ͷ�>��߻l9.�n��#R L[�,
Q��>7����hu�#q�\�T�����L�H65*x���*P@����G��^���N�Ӽ����(�E&�}��^@�ş��˘`��:��8��E�+?�1���Wyys!8oP������C�!|��ȽK/1���^9�!sW
<) t�L���$����'F}qK��vQu]�~
>+�C��v!ד��������wZs��o�cfb�B�o�bM]ww�S��ݞ=q.�z���z׉�W����ø����K O�����6�r}��w����3n
��bAb�2n�Y��&s�A�d��m�B� @�g��w��Y*���xn��k��զSru]&�<i"4�u�kƳ�r�H�����7E�u��3���f�
����g?�x�3�{�N�Ô�o-��޽�0l9���1�tZ0���ӂE�2�X��$��Sd�uš��X6php͈-=��$�nP�Έ�^�
:�JN&	!k9�f,Lh�����NC(:k��қ�F_�6G�̏����(�9�Hs",Z3�����������2�ӀU �Ѧ�_d�#�<2+���s�!tv���~rd�;�	�^���t�ir���'Qu�H��Z�����Ԙ��f# ���Zd��.P�pY��։�>
���.|�U�T����o���`P��%�h���ܣ����q�D���;g����ۦ��._3�?���4�S{�gW��Um�W��Wn��=UP��$�Q���J&
V�YflR���]�C�-y��c|���K�h��}��}�*i��U��A.��;�?}q����CN�Q%�{yIY{���v�j�H�"�y���y�bfQ^���T�hQN��MV�123Gmu�~�y�{p�y�����3tpȬ�$>Xz�Z�͈���iQW��8��m-�L��D���4Ն��DC�����0s�{O���D �nk�ĝ��CN�lq����� bקއp���B�S�<�E���]���
�1|�5�#W�><.D�B����KZmw�()*� ��t]��@�W���U9�-���O�UO}/ijp��.�l��(3�h�Kjq��֕i�!�6����yב!x��[2|�ҍ���3�%p�DȜ=5��ʊB��@�9��A�Ĝ��o�H����K;��&5�2�1��f����*�Sb�${ptM����Pg"LĔV�����<�0D�۱zU.z�W��C�!Pu�.>�@%���f��g~��9�!ԁ5O���ƛb���]ʝ���[>�]Yo���$ܽ0��V�eq�B�B�]v��?�*�|?�8W[�2�'�Cvk�°Cc�r�#��v�R+qA�Al�ç��U��־�E@���"��'|(Ə���c���?�NqrZ��FMb�~�-�F�����֛y<LT��N�)��nr��Z(vEٌE��9�Z����I#��.e#5�