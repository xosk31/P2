XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����R�.�w�<!�AK*�a5�4�v�	�9x*E&)FW��B5���[�����R��J�eY(jY�\6蒞K�-���r�J~���❁�B|�8j��'��Uxvu[�>{��1[n�g���߰�gs��z� ��V������謦臍eBX�![t���LVn����nE0�H�l�k7��յ�Hn�Q�:M�J�S�F��y��[��1|6�(	�Bڧ0���>0fC�?��Z!���o攓 j�<g�:[�݇.����g"n���-ā����M�_V��XC!9��� 킹rr/j��7��R��Y�k��)\��B�d(�M�.�!R�*��B�ßC����*�(wj�x��fWB���W&�E�`t��7�l9O�J�/_/3b*9)mx�Ra���,���w���ShVF�p<ơKLƳ��	cqIV)qx����Z�U���h�~��8��^�*K�5�y�M�E
m����;VE}����Р*���⬅�������.��`� �ŕ���Y\H_U�kNH5?��<��fW�����s�\��l���z�*���vT�{��7��m~��xulM�@W��3��<O)Z�5}y�z����66����=Ô�҃��rt�Fz�
"��<��4�&g��iɈ�����v�y�A�[��o��n��̡`��U���5�`no�'n�LC�d�d+���/�h%��/q�? �l��T�	� �!�D���3�4�$��h(,]d�a�kGWXlxVHYEB    2fbb     b70���p�U�.k�̔�¶�v��e���@DL"�%7����n���9� ˯�tGS
���*�6��0l|���+�-hp	���\&[��m���hʦ��s۔���?C�������ش�F~���FЋ�G��j��O�� 
F���>ߤ1����b�[O}�m�C��x ����-��,l^���أ9rr�$ɣ{��x8ݞ%�6)��*��j
�W�	k7�����sf�RI.���2�H��f4]�-�C@��y`�*n&�A)aHJ�P#^�� ���*��e��9�Kկ ���
����}�P�0���dD���r�A)v���8	e�0������5nsfa�TʩL�y{�`<�^'�yn_�k�Թ�xڸ���[�׉��Q�jE�vBu�!DH�3ϳڸ���1�R|Xդ��*{��E�&�;��t��N�{���[_��퐬+h����-�S� 7�j����#������@�5� �HI�0��Rf�l�T�=Cٸ�6�rݣ��r�}/d�g��F���c���G�܏�T�7DB�v��y	1M3H�BU��ݽ�]�W`���Eϸ^�?�������v�\kѲa�̹��^�K}Ҡ/-�,��Ii!��y?�r7b�Ӷ%�_��9Ӟ�禦�.�Zg*hO�~?����z�ȳ\��O?�J�	 w�M)`ݍŵ�T��)��ʌ������n@���l�Q��©��T4��0.�@�+�m�#���Q1@�/E�ޏ^�C�B͵(؞(� ���@�,�J�-@;XN�XiT.����M]z�C^���=d񒉄?p�k��i%��x� i��}���N��J�lx�M��X��0�A~�0����*VgC5��Z6��*[g_�yb�*�e�A��x���˛��v�fr��#�?��Yff�'ۇ7/�d��tD�u)�4�:q��#���`���'��T���٥83��]`��d��x�/��m�D�a3Z��@��T>�������z�ʞ��L�bID���\�>�h��$!�|��7��HkD��`�SM0D.�� ���H�OkɆoY�@9�Hn��q	��(�jw�	>��常�JZΟ(����<�����x$CXy-p�D8�G��=nt!�u$	a�<|�fFخϹƅ�9 ��(Y���cu��A~f�>Ak�q��P�D���!�y�����{�����<͑�$#�S�z�hzT*?9]����r ����).Ϧb�P�X�4�R�6��:%2�����n��V۴�;[��r����C�?­��Σ���n/����g�%�n �<7wc����ѷЗf��N�tɋ<�%ճ���_
/F��[��˷��/�'�r*���-z,�']��!����d��rQ�)��0�?���R�*ݍ��+�'A}����7Az`;
���������we L �zF�6b��3���`��G�KZ�
�LL���'n�[L(	ԁ%�y���\��!�n�̋������b������#�K�:kBP�
�������6��nt�Q!�X�$���]ЕN6U��#�[�	��n{�4�d�5��Qd�jYK��i��d�&oɕ�cPW ���T�	]v���E�F���!��*g��@��wvg��8B�򉴭h�aK%e��;{%���l���('>�V'��Qujh�˟B�TD˿���Y����8�����]>$��΍�~���j�~��?A���X	)\�{�@>��e�U]���e�Ck�q �I�T��&�д.0z��UNNe����W�g$�{l@�^ҹ��ZS�0iI&X�#3n�������"�ĕ��&\6j_l��K��L��1�c��s(cgB�|������ycM�?�:�ka���t��0���dᢟ���:'���bw@�o���h��&y�u4q��/���̒}����1�0���������Z;s��˖jZ"����Հt����	7�^iti;Q�pmd{����&�N�Ή��EfܞG��Q��|�k���Q�}���#Bd��^,%�#��6^jH8�w���R� 'G��Y;o�x��e�ݷI6�ҡ�Y��k:��ˀ���7��1�G�?��I��3�9�p�������f �'���M���,�,f�8)�P�Hg �`�S|*��+�LR{7�H�ǅ4k?�� �Z�&��$��kQ)R������5Z�3!u�eE�<�k�P��b�F�'��>�D���[�ӂlW���	��7Mm��� �� _�g�j �2[%�����U�b����Xh8��J��_rں�6X���z�R�Ǽra�
r,�K����jF��\_)��_�qW�jA�^�͗F���>�嫲a�leX7���do㒅���v��Btrq߈+����J�f/,�.�Ԋ8���J)�zTbx��������պe�.�pD�F�c(Y��T�הwX���7��'�.��f�G�� �MRB�����_�Ԛ���2�8�A�e�#��ps�m�|���礩ry�,��s�ϕ_�>�M����(bY��ݑN�⋔$$g�|�����zfK�a��]��E�����(5�بs�ԙmwSѮ"%���.�I��Ҝ���@�$$[x�S�>0~ɰ:���X�?����0��p�J�*w=Q�dE��#���������[���'e��2�A��_X^W4��������x'��Sٿ���v�I�-���M;ƵkB
q��3���p9���_��a�|3�$������=���u�"h(�3�����&��6i�@b:�&��5;��z~��&Đ؋�Ort���j�}{:H������N�c��T���Q$�q
����l2F���3���nL3v