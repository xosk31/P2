XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���A)�e���x�vň���=�l�����|��(Hk�_)�Z\d����Ku��눤�M���:�:]z�=*l���' �A�x���dS�-�~{36a�*����}j�J�H���9=�hӼ��`F�Q�/��X:�z|�es���0��>f�{�!�E7���4!a��{�`����O%�($ͮ�Tc��R�6�Kp�$������)�w��A2��Do`�i}��F��Ň��A��Y��M��sR��
���5��H�9R�	&��d`1�U�֥e��?�d��k�V}��a��HO��l�o���Kbo�pZQP� ���Ɂ�-���v����y�����ٮaCSU{	s��%8��~������~/Q�65Lt�z�ҙGx:�M�ɩ6���w4���
��$�t��m'*?'H����wJ�U�H>�p��@�y�p)C4�k!����uvh��ժ��<&��]ק�6��#�/��n���!���`0ͅ�z܇����ذ�_��?5��t	it8��$}�p��a�"r�k��Ө�*^�M�?ĽϸP�6.~�VT�R�(V����qܪ{�H<�����GoHǇ9�o���Pt��l#̝�1��͟���}8�C_:1!���>Q����N]I��Cy,��t�Q�!�5|����ʒ:cr��踦����~Xx�̆��V�xL^�?)��C�T����?���)y5��80�d謇Øi6��U�m�����q}#����ᤤXlxVHYEB    761e    1770FU���=�������	oě~v����D�#/6�{F*��_����/��o��÷l�?&�-��cqT=�Q@B�����b�w�`�G?��c�a�ɨ72��`�U��ӗ�ٯ�'�:N�DC@�uc}|��B�_��3��&�u�8Ѵ;KO�%kSŭb���V�r�[�V�� �"lqi��Ùl�G*��R-�.�*9���
0���֞N�")���z�B����%���$�7� ��?��e��Twq;�<Q'����)��n��M��p�Q�;�\���y�N��7"7���߷�|=w��A����V��F�ݟ��M%��.9�Pp"����""��PO;M���|lc��Fw�dp�AC s��b��F�%g�*�7��IC����*��Ƣ� =��h���l3�ճ�{�RJ�i)3Ԙ�*���tlO�Pu�]�� =:��|/�s�L\}�X1XX	 �	Ѩ�'|1~���:�u(��G"@ട��s�������N�����5���)���0W� �w|�ٮ�=��1�),	~cp3�˧T� |���1�C�usbAY�(F������s��a��Ul����iQp�,��h�q���{T�B�"��X�� i_Ǥ	b�`�<i2e�x?ݖb���^���Bo��a;�����eV>.��}T.O�僕O2�JGiAȍ�����c�j�2��Z <��ڂ=�R�?�s"�~��*��Y��<U��Hr�=N|U�9�*�����mϔ3��+h�T�0��z9tQ>��LjƏ���]0�}����;P#1�*�i�_Ӽ�QV�?6���4����~��_���X�E:��d�:R�e`�A����a��|��n��?��uGIeYo��$+�9���B�g�g~�>��m!j���k���T��� ��ܳk�0[OR>G8�B��ͬm���=�=78�
K�;ӄ��~�u�V�KP0�!9~�9^�{{���)2EN��g�96�<�Idr^D8�݉�G��(6�#S��4qȳ�7���?Q���	T��Qrh�+�|�Z3nM��%t��}VarE�5�;�پYLu���z@Ö��5�8�1�'u}�m0��v�./�u����rw�\�<�C�����p�KQׇB���پHc�L�q4I� ���n�;T\?Uq���
M��C�U^x�L���L�ȕǸK
]�
�7/"zNa�jBE��\<�
?�s�JS����>��5�r$�G�ڲE}���J�6![���ݥ�zN�@�#�9x7���)X<$�]X�3+���o�yGAah����ޕ�8����_8DE/�:���>5` �����f�@j�o��},��5��pfx���~�p��J�pn�E$�9?:���I�G7�/�\���d��1"q����@�|k�]"�:3*�`��f�O���)��8Xԑ��J��xf|�/7�!�Z6��k�:S�b�|:�; �5��a�6Z�kD��-S�M�c�����F}ms�]L��HE�3�!�F��OI�U?N0���e�%��C�9*0I�R4 rB{[j�V\]�[SI !���7�[w�!pU�d�'�f@~`�{�WcK���	+ʻ��:� ��aU�&��.����c�q����"�wc�uh��1Ħ���+ػ��KⲎ/�ш6
�=ιs��%��9߁�|��2*�ǅ�}}��c~W�<[�g_ʙ+m����z�A��`��$5�0��K��g���;x&ek��ς 3[��	pμ��%���:��&����!�`K)��폪�A�8J�<���]�$����^��ZijI�!E�)������/R;��h�>�!Mq��REF�`������U5����f4d�2����#�ݒt��0N��i�ֽ��6	+��TĊ����"צ�e$nzb.�e<��{��f�w����M�rq��C�)2����Od;~ٵ�C6"���\Im�e�|D$bؼ/�����K'�}p�~���}��W_E/Gp)�j#'�
�?Q�������6j'��17��M���W	v�᎓Ml�MT[|e� �q*"%��!�����ѧ��Ӿ���/ٕ'��d�W�ho忝<m0A�c��6Śv��=
^�"�T��q�ڵ�Н�L��/^A�����ݗ�P&�>��������0S� ����ƚN�d w<\�.B;p��Hz��Y�Èf^���k�ܒ� ;���ߦ��6�A+`�g���g�F{LC׶WT�j�S޺'�N�i�t��o�qɠp��`�"��]%ځ罙!��Q�~ɜ2�?���:�����C������ef��ko��%ع⋰4!�͆\H��j��O�9�	�thP��ڂ����G)��_�x����lJ��i�:�˜�*�@L:����`�z�1-�J��OQ���|��༉���������P�wƑG�|k¡೧1����i(Ƒ����wg�ņ3":+ᵕ�Xk� _"_λ:FCGQk^�m0�N>�#Z�Y�Ҩ�N��'0��p�M�A-`��s��Tx�F�p��d�$��I�0ɓ�ӳ�'��A�P���^.�ZG	�17X�|�����|��+������d��H�졿c�g���mމGzDk��N���CV�^��i�Q$�M={��`d� Y$�p�����2�YO.�����Փ�.�x��I���Y��A��Qы ��?�K.�yg��`��(x3��+�R}�F�����)��dDw��O����v��v�o��&�,���V�"�|*ںy#�W�e�>X��)_ߧ���[z!���華ǰt)�"n-6hm�-y՗�%��L��t	��?|���m������� 40�`�x���kFT�	�Δ���|��Q���d�D�F2݄��-	^�?�=qD��8-8H��̈�t}�ɜ!N����~I��k��-�ђO��cB�ҟɔa�E�	�>�"������M�I�S=)�ȵL�-]���`�_.�B���ƵL�$"��іY��hI�PI[�ɐ�Wg���-o��N�� �m����y�MJ� ;�i�N��2��$�� /���l�0{d��� ����ź�NPsAZ�M��&F�M���8����/Q�a��t�����x��z�d�C�`�&}�8���k�3���ш)f�uY��%`��on�.3`�쨖fC]Wxi��p��	�Jb}��x[|x�.~��GK��0f�2�1G�ldP���Q�
Xs/�((4�ۛ��Mv\����~֭��JGWN��P�X�E	�	*�Q�]_��%P	�q̘�H��U��QT!�[AN�,�[��k�,�`C�:����|`�R�޵l �U(O�x�	�k4�Ө�M�o`cF�[��X��s�L?�~P�niPN_c���6=T�p���� ���d�9;�����|V��u�M�MP���lH �+z���ɽ��Mf�D��dMS&�3��+���gɟ�����[�A�ST>�nS�l}����8���s�+I2�'y9k �����g�@;��ۛA��|�w��?Kג����\�ǦΊ���ԛ��f�skxt)�h;F�6�DEyrM@J���f�I��h��O���:ƀMp��L���0 kO����%baaz��ة��Ƨ��Z,�]ȟD�����m�J߉;�;Rpd��GV:�yPpTסӶ-�œ���b�s�ר�a��s����J,���E�2�Q1�~���R����-�{�� qXTӠ�+rCBѭ��������$ru��ܝl~��^��ч^H��J ��q�,��1ꋭ���!Ē�j�9��+�B#��TϰO:2��.�l������^,=_,#��[~�.�����-���it���0Z�$��B����+��t�_�dۜ�\�������5~(q�)�Wv^��{���U��T�c	�s)b������l���~/P�
�@=�[�A�=��ț b����K� �<�8@�!�*�+=�L��j��j�߁�7nt|������� ����`�e�HR�����a��Zw>ݸ�>M�2�����"Ќ�v�4��O����x[T+P����Q[N ^�����ej�|)<7�w��I�d�xM��Y��ۈ|�Qq؊�6A2�\��R�W<8��v�O C_ƒ�u���)
���]�/\������V�S�k`�n��'rH�*K)y�Fz:��B3�+D��$���B�Єt�ӠfC'��`_���v��<��p��Jx�c���{ m
=�+�|���5�f-m��Hkz*
�����k�E�>�����+�G̠�:�:f<�!&s���4�66�C��X!z��<ig�#�G�=2��o
��,�<6x�C�"�n��F/d��h72�9:W,����.� �$�k�ʅ���2��Q�ֻ1��g���&PL��/�|_����uBP��R�*�Ϸ�h{ Y�R��a՟3�4yv��Z�i�b����[ȓl��ɺ2�������]kz�-o�9O�*awj}��>2��2d�高�A|�!!wng�e���(�O��C��:�P5S�b��])ڱ�T���&\�leV6IX7c�Ϋ�l�KsP�]�L_�u�_�� o&E;'-��"���|�i��^(AT[z1�����w%�,Q��<i[��[�f4V��l���&��l����n�+��{=�;�Ϊ�a5i>G�=w�-�&�VX��\Y��6C��Z�K��
����k�;��EŐ��c��nln�wV�lg`7�Q���p6&~z(��A�x}a+Q��h� tų{�l3{N����1�����Z�Ҷ�,���G���A��/�TrGג��TEO6I��9&Z��:#�=3F�>�ˣx����N���/c�4���3���4�9�4G�H���nDu��?�ՔV*��	�Ge3��kW';������P#��x��`i`���9ݬKEWX-Ǝ?	(T`BM#�NBG�[Jۻcƈ���bh��S[U�ry�GՔ&��Nvt6t#����)tRe0ҞBrX����Q��S�D��7\2P\3��=]O�
���}5V�&������!�\׊�ZE��+~x�� �۪迨��	Y�b��-�\��Ie�
�t��8|�{U�G�ֈ��,c�	��e�67�+���<|��[b�=;ȫ[�P�@�2�r����Q��O��"��	L���/��	ߝI\�ᤜDK��o�� W#����0��Ġ6�x׷��*=��0%�'�	��7n�-�K��� j��Y��B61bK��?��\r<2I���T��<�t?wȘ֠��5��!�������8;S�	Bi�K]]V����.�N�Y��Bg�`�3�r:�Iv K�̿n�t8s��0tnP����-7��7���͗���� ݵ�7j�'�64�&IF ��X���S!���^�&"D�}Ŗ
9I��)���;�Z!t��x����aR���j��J�K�����V/Z�&jϛX��[�M��+d4>�`�����P�&�2G:N������Jc���9��Yp�U�/BD����N�G��`��4�_�	�s/S]J�\�����	P	01��N<J�������<s��W%*0��8�+�a*���cl���ksY[�+~8h&fz/7]�:����\On�a�rs>M�_d�K9p�	�"���`��չl'�t�C?9.� �5����I�$t<�������j�G�u�M����m�A��X����*N��"8��PŤ��0���bA|N��~'����y��m#R�Q����*�ט-��&�ׁ���%�sTn�'1��d(.����T��3����OhD�
��j?�����E����Ӟ�h:����yX�e