XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��pfyduj	<��Ff�,�U�o;Ԙ�Sg�F��c�x�0�l^�;&����(/�B3�r�)
��Ja.�,���9�F�4r�ds60�;����&�g2��U��\���E�������Gs�⍯�Jh �]bc^�o;vr�u�.�y�eصk��ZFz���:��-��,-܎�>op\_r�y,	�!�I�8��O���Xa��sҞ���́�� *����������*�?�yH��c��3	H�w�S�`�0h��(���m�[,��}=�$�_�2ΐ?�veW���É��9�6� ��ngEǟuLQ����-�O^�`�!Rz<(9Bc�됒��4�ʸ���/J����!�s��ߍ�5H�Sa��M��a���<#l�]�[�����?�P�4;���&��Yd�$QnI`;�?�&(����^��MP� S���$g%�b��Q���8�=U1e.�jaYS+'r}70�rd�|��:X�-)��SY���4���(��c�i�F�^~M<��k�/D�xQ�w4�ϙYȖ#Pm�>6�*5���N��=}�?C����l[q��u��Q��*�(�&&
� S��*�q����V0�Ʋ�9���+tc��T53�E�[�Kv�݇;^R��rL8��i�wqUԜ!!�V��	�)�S��!��5�� ���)����1��V���5 d�
@X �W��Je
{b��"W�BS�qr�0��d����x�c4�f�{�����@�yeXlxVHYEB    8990    1bc0y��yr4R�w��r��M����i�q��n6�����y����k|r�j
��L�z}�?i�Uc���{������B�4Ee<�K�R�ɟJ�y�
���v"تC�:%�8)��̠N���L��&􉼦.kr�a�,��o=�ߐ��¤%��!��,����Ɣ���(��,��$�}n"樽�$U�)cl�n���9� �]�ɠ����#:�a	��H������oS&|W�^�!Q���s�t�A묃���߾�9 q���8#� �N���!�S�����S�l3�vc�d������n�*��o=�G  e�ަ�������}õ�l�,y�����y9�,]�D��y��癠�����˔�k�����ws׿b����M�Һ��iV9ʨ7	`�[k��Z%J��1�^�Dy���Y$�`���,Y,��9}����VA���!��:�+�-NxxP\hH���u-z�\�m	#iI�E��5��x��BS}��S�3�b�r��i���#�%]d��E�<ԫ7���o���0��LyA�H��F��.���
q<=(�ܲ��FL�(����M*d�ɻ����S���D��f��խ��ډs@�݄�]:94���D��\�y0�=�#�ˠ�����8��X��켳��>�Qy�8��?�Tj��P8��Bӄ�aUL-�������;Ռ���n������s_g-R>�v:-ń�aאK;��g�֖�3Ai0�s�
ᝯ�Z���̇夬�;��5�C���M�`e�� y���C���	�Ӎ�q��a�03R�7���ߞ�2�x%�~����EaE$o%\�	$�xܸ�~�4�L���Ĉ�!��6e~��'�L�I�x�ܡl�zt�5=2�V���)�1�1��y����#\�@Zq�����e���P��i�pAk�C�ի��D������lM� ���8׃�a��$/e�x�!Ki�KCa]R!V@v���W���Q�M��|6x�G��3X�&�����ǯ4X�#�0��Kz��o��P���EoM-�JbɎ���ܔaq�i#�󈚠�� �;1��,/�1�0�f��n��=�ڒ��8g&���'o�L?�4@G+l�P׆!9��	��/�\@����pc�X�2b��{��̸0����ܘ�<��r���o����mW���X����1�Ժp�"%�>�h/ �R("4�ȕׅ�5�F�ct2b]u��ʀ,|TJ�n@E�ZP�6|�ri�����F��Ul"o����}3�JV�.�!!:�Y�ete�3pw&Fn�_3u�7�1��nMӽ��n-t�pgZp~�ҁE}��.�����֧��ް���Nt�!�u���OC�������묦G_f��\�#Y����$��_�'�~>���&Q0���uEU�p�
o�1��Y��+f���{���Wƃ���]9ѕ��nת��v�l�+�g���[T���(y��c�	�i�}b��j|9��u(�1���Ę^�]#Xڝ�:�x�m�~�ڛ�i7|�eNx�|�'!%x�t���(�Jɛ�f���\�����:��;�]眺��� �!:w�wÃ�?ɧI)v�/�V� ���M^���1;�Z�E��t���|[2*�7�]�]S	A7':�]j[�[��۾d(m,]�G��ײj����u�.0�	YV|.jn��Q��8��,���(5�Q̛&;v-�|����L����J�2>�4�y�,w )%1<d�[�4"G���@� ?�����E#�}��C� #i�̝�'v�W�2V3�l�M�p
�Pl����b�:��j�B���C��u#JJ�yʈug���倂�|�d�;Ɛ��4k����� ����c���UdqPV(9v�8T�;G&Q�G(�p$�ܿAm1*����fc�����p��aF_�Z���}���b	���v�3rշ��x��>d�.�	`-�g���f�9;A!UJ{ԡZ��䱎�]�C�(:+ aM$��0��[����������%�H�٩��snǼM�����G�nՒ���~���ѽ(�F-{�1Q�{�,�A�w�_c�s�����Y²���c8Z��Q�S��R�.�岨����6?�עSؗ��Rf|?n��*���k8q��0�.�f���1��q���hl��^�M��j��a��qJ����bJ���u�����]������}�:���C��<9��q�M�б`m@U�y���$>�uG��_�I��T<Y�/^��Y��9�A���B}w.�Q���J�<�ݥ*��r앭�>��q�L�t��D���>A;�O�_��9�>~zҎO)3~�n��y
�>����О%ix�G�^G���d��0�53�V���̶疭��JxK-�+O ��z���hh� 0V���y�~�4(M���<��p"�&�E��� A�#��Fu�ge������k���b`�J��a��՞<n�%!h��!���Vf��`)��>fj�*�R���=�6�$
��QTSQ*����zZ׈�+�)'�~�Ҭ��+(�ه#��~���
�Ā�߻��ZT�z-j��v=2��<]�	>_�d�Z�S�����Tk�
�N�~1y�����W�_9x������$��?�>�FɃ�-F�xC�0���;4�]�mST?u�d��C�$$����M>�QqM��\���<�j�IB�t6�9�������$|�J��Q��ڭ� ������s�n:ʞ]�\���?�Tn׃�/^�V�]�3`6��k4R��1M����MF|���=��SH�ĩ�N�� ����T}�!�Y���yL+��8$��QC���QG�ޭ�:�"��G-d�,��/lC���<�p��|���
����e�)Vu��>����Hy����	��@F�<��W��#U����6���~�1kژh+��y�
$��I��"H����`F�4�^��@,��ZTd��I`J�����h,U�j�f A�1����~�<��N@�d����:�]j3�;��/����n.m-�$)��k� 'b$��A7�t��j覘x���)'�j'5��	�7����\���H�����)܁u���(��q��k6�13��=4�y�"�'�_*�F�W,�l�����K��`�ᚒN���@Y���9����L䏾,������С�Gݟ��(q@S���%��ڙ� ��I��)*��N�;��7$߃���4HQF���x�>#oE�`)V�o�E�>{��p�7u�'�:Q2����h�A���o�����;�+�?�O���ܿ^ʄP-���)u��c
'�KR�ag`�)]�v&��#_P�@��������t��kE��	���cY�d�e���h2�-��U�u9��Eo�bK�ߥl`�VŌw篻��G�J��0V� |:�
NA|�[^��f�F��_
i���kD�LWn�V�x��;Z�(zu��s
����l;yRP4�d9	�L-ŒK�eX�oɆ�RԬ��Xh����T�!�۞�(y�!%����ri�P��c��ۨ��_�I
�3��*�� +�%�$��(;�JG%�E|�♤_�xB��Ȳx�D���=V���φ��G��0ז@�F ;yj΢�ͫ��S0���Ǩ�S��9%%ε�� SC	���v�p9s��>[������#�iy��Ʋ���q���V;� �ty�6�:wLWx�N�2����������r{Ъ�;'6�κ�*��&�҉6�ȹ������t���k�����p�T�]��(L`�7���)���CWn+��q0RY��ꐴI�I�jA�^�W~��}�o����͗�,{�̻&�0�P�`��Z���}��367�bL�� ��\��A� ��Ĩ�Y�߻�r;;<]�Sg�I�u�|�O2�l���n뮛�`�:�o��Ab<h��p�t����Ͳmj:?E���2���b���ғg4%�	�_2����!��Hl3uL��4�v���W��G���R�ǯ�:�'P�����>�B���pNzS������[���&��[V���'n|��3��g�����
�-�Rb���r�y�������#DZٽ�_�u�.�뀑�.~<q��&D�9C�1���ͬcG�%�1:eC�~�E�@%_ �?���/i�<�GL�y�#۵�ԶA�X�����q��#�czV}��yS��li��`lݳ]ڜ�
t{��~
������`�M�V^]ݚOu纝c��=�X�N����`�CZϙ���i�䛆/�8�gr�{���u�D�̓��\�x�c&7���m9�� {��ᾅm�V���bȫ>v�PF&)��*�r�s�?���n�f ���y�;K�'k}>I=�F�wT�,}\� x�|T�U�B>`f�����;Y-���*�A�u4�x�ct\�§[M�������[�	m�7�Y�Ӗ��z�Z�׉�'jr�ows��la|e�?�MV)��0
Ҕ����l�Ęٲ5$�,��ׇ��ڿ���ZB5"����S�ve�̽W�������S�E��:��v��1�Y.$�vT<n��U� %	%��+�(jv�">l�4LOw�ƹ�t��Թ��^V�X�cH7���w0_�b�+ ��xIPn��m��UTn{�;�t,Fق�ْ���8���vքJ����.3�*K�	U�]6�Y}�u~��`�q�P�$�Sr=<����8����g�j�BYڑ�����Y�ڂrʨb8��c���[��7O�Ў��l?���g��t��R@��}WCU�O�=�Dad��� h�;	���L#�E�/K�WN��M���J�ic1�, 6@�8uM��=�xm]mS��G���:�_����^޳�H�E��(.�K���	��~̟�"����v\<�~f�8��JH��IT<��UP�uvZ�6^}�xEJ�-��Z+�u�2�*��J���|	Y�nW�~}CrL�	�߭�h�S��Y���}�{��#��ZQ~{F�C�Q��ٳ��)���'AC�u�Z���F�,Ò�M[�-�!���A�}��*Iim�a:t��~�x���r�Җ�6��u�#I��˓QV)o5x$e�u��_�Af�҃P�kD\������~�o:�@8т�����-yj�ζ&^EL��e���yǾO'S�e���EF�nA���'�!��YL�[a�3Iw��bRC��~���c.}!�r�n$h$�Z.���n��VNL*�#���+����w7�H��CU���x���F(�E��� ��7��079c��F�ʹ�,�D��
�>�gN��2�->�';��60,�x���K���fh$����K�������,g�ϐ��a��Lu� ���b%��91�ia/C�>����������W0����\�F��~�X��Ś�o*�
B�L	z t���4m1n(�|��,c�j����ȫ~7�b�Irf�9�X�s묙�I��`�~ﻣ�����!	T	�U��LƲ%t�%Ex���52�5|$��$�HjxKj�rl���d�[�1܀�͔/>��k���	y]�s�i�Ikԉ[�]�����' �Q%�F��^M7R[!4q�Y��:�(#���.�o}�[�Ve4O<Ĵ�V�v�����[��y�Mx����JuD�=ڼ�f8;fF;MM���>p{������Pi�د�"8��^�K���<C���|ɯ)�i�R$��p�y.��Xo%C��bM�|�m �Q�m�lɘ��E�ʩ�a)����H�B�"T�p8��Ѧn#��:,4�E��D��2 1��"���{�|!�y�ȟ�0��t�=K�hK$� 9#�!�NMh_^}P�<�|i�;��ԩ^|w�#l�N!e��P_>~ѭ� e��R60�<${��/�a�O@���}�ys1O;{�n駋�0d,P�fxn'��Iq)���ދ��h���71��
So���|��f$x���W�*4^Y'��`�<Yd\�+�&���	ral�Hm����Xu�ji\��.�u��ą�����̶h%����)�իT��%�\��#���/	�k��=�b��>�8��iwP����Xy���l��4�:��c�%/ګ����y�U�-*�8�����o&`>�ăr���	�����{Ɍn���rj� ����E����g�<���$�s��z{I��4�,���C�/�q��^�f�_���%/���D�L���&�;��10$��O��֠8� ����
T��� �bf9'�9�b	�~�+�]�9� $�-�f�����0��V�n&=a]�'w�_��C�qbz�Mym�����쬝Q�S�<72��݋��Q�S�6���[�sྣR��<���=-0���z�޸�������9M	��n����݈Gv�]��4�}���5^7}H�E裄R�Z}��l.p{]����M�����f��������R�����D���J�sRcU9$�>�tA�V�H�|��e����ڶ��j�y����)x)��qa�)�[�6�L���˧�-��Mi��g��W�7/�ĸ������j
���E2Ft�`�����d�V/�ۢ��&�fK`�xn�oc��@���w�-�C9�tO�����D�	�!8�cE��� ���;��1��*���̴���0J���mo��簉��D"�_\5هq�'�k���y�/����&�@d6�,F�Ns�	@�o���@����E,�D|���d�U�������`��b�����.� �i����KMR�x��1> ]�Pu��e��Kgؓv�N��h4R{GF�e/s=�����zj
�J����'O�ĳ]�J׼~y�`G�����U~3�62�ᅝ�D� �]_�V�؎7�oĲ��ӳh�������-���,l�ư��F;�.�5�R���E�aG��b`���&O��s�@�7�?��-���k<Qt�c�J����K'��̗