XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��7�`~���B�	0.f@����|�	/}��\!�GK�㲺d�sK�RX!wCe�b�M�������:��\:��UUY�"B�ؓV�[�>�)��/��\��N*�N��P~�&��(H�Έ�0�k�'�f�e~��
*@�L�l�����֚,�Vi�mH$��Ȋ� җ�1+��BBB��[���F�W��#}�\!Á��]�X�B>���>^}�6����B����PP���Y��Bk�����[ �f0�Ԅ�dx)��w����}}�1P�0$e����+��^���bގG�>$?A�
/;8�� ^h�+��ԫ��
���p�řнY��ɇ���
�e��)���	~��ݢ�nzW��$Z���!����Jp��K�'���2�i��6^Д��O]'+�L(�p>����}�j�f%��C
�_�sk��|�=l�ɢ8�= bD�I��sd{��g��t�,.����b�Ec0K�������yI��8�u X9�7O;���I�����1����1u]�jh@"J_�O�?X�\9a2AH�K�9�'"
�	�����%پ�TfTz:��+��0%	�FU����{�ccr��yA����wIE�Z<����u�*�pJ".�?"*	���6K=�;��5!��J�u��e9}#���D|):5��ы�鵸�:6i����}1W���]�t��F��:q~ �q(���6�����ٗ��Μ�w���ݰ>��醅���ӓ�s6_M^ �<Lˇ�&�QXlxVHYEB    fa00    2030QI���oO��+��
����
}�'������;[���� t������mRd=��<�4���iu���k���,��>�T����[�yo��GR]gK}��4�g��@�f�W���g�<�!��Υ�WLZ��6�X:y�����	�H��9dR+vb���\&"O�b}���hG
R�{�2A���+9"\O��4O� *��13�g�������<�]��\�C�\ePl�\��M�O�2y�( yd#(ޣW��UsR7;G�AB�Q;oT�L1鈠ѽ�0!J�C�$��W�b+\FUH�{-P����I������<c$t�&p"!y��=I�uH��3 �/�W�a����SN��Р��V��B	��yu������'ہ�Ő�n^��TEC�GP�͔
������~FXB�u��/A*P��L��ؔ�'�dw�ū�;��=�G�M��7�'�Ƿ�&w3��<���!.Ð>�xgI$�1k��uR�Y�.�{���l�ʠ�)����V�!��M���T�.�d8�M�jt+��'Ar�U��6��:�KW#¯��h��O�p�:0Wqy�*J-�}��[���(D�CRCX�mT�?jl.��>R�J����,�����t�[[�waF=��k3��",�$����5��p�y�bZ�r���,����7ܴyHY���������1c��W���tl�Jj�!<��ò�a� �� ���8%/�v�jrW���h��N�d2����c2��i1�突qG���ۂ��K�Nk��S���19)d��&�1�*�I%�B��jق�3�(G �	3��uԕ��ZV����'����u+�{N�<�R�Ƌ�6c�$K�*}����"��ݰJ�$�����k3��cɿ�3�}uH9��}J"^d-B�lt��l"�f
�!�fk���8d�L��4GtN4�NA�.�\�� �j�Bc7�2��,�X�3Q�O5C'ÉA�^8�6w��l��?�Z;�����Б�D�nF�P�����mϠ�뎦Fw��N�wqu����G&+�G({Q(���uYKo�]j�[dhk�E��c���ϗt��2��S��������IOKj������Z8�<O��<��"�Z��!S �	������%�;Ap�Kq��":�0�A7X���L-��;��Y���ċW>ڱ�����/����ㅡ	�g�A+&/B9�L�=��I�٬嬔��j��1<��i`Ģ�&��Aw�χR1Z�֡�mtX���!��ﱑ|o�vZd(D���E�
����M�3��Z����*��J�Il����I�3�V�~]6��D�9j�`�9��`�j�}K�ĺc���(C��v�0�}�ȥWGߴ�� ����M0dE��E��-��=�����~����S���Li�	[��p{{���hȮ=�̲\������B���/J}V�{�A+�3.~�\-�]����y̟���#�צ����79�К!+�^�o:ϴキ�C Md4NJ}k�S�'}�ǘ��#�;�% \��o���^���~�����Zt�	��«�S�3���
��9�g�T����A�y}��O�<��5
g֬�����W�j�o�ּS)�4�dnJ6�z�S��E��X��B���	|��S�mӺs/u#u�Q�>6���u7�+B�'�����`~#x�(��M^���u�µe�����;,iW-�*Y�ʋĀ�°2��k��˻	X���E���Sy�ut��Ĉ�Pr���Y�q\��xR,�����bZdq��iZ��<��c���C��JVhFFYB�CI=��*��hd����@����c v��Ek�)��3���� ��:���8J��K!:yo�3瓥�}��ע�Z-�x�,���I��U=�t�pZ�O��cE�hsr�сm�qW��W���Tٗ���2F��MSv,j���΁:d�9]���ݼ*�V���a ��#���g{��>3�X��Ap��=��`�W�)p/i��Y�r��݇[�C�d�5u����(�������NAvx]L�]�<��E�� ܠ���5�I!��:e5}]A�ğ�NA�kXo�*��;R���#)7-��ׄ
�}0�i��&�"[����l�o9��Κ�(�i�����()^ѵ"N7��J���´$d.��v��>N����)���֓���Z�����TB*b�Y�ðR"+N�/�#�	���\���,�{�R-�rU� ���II$8M�8�V��z�FL�:Iい�t�zr��hTf*ܰ�ڳ�a�)�ӈr����)v`ќ�e��_&��v�ϡ�z<#;'�Vj�ɞ�"�+�n��zC�/0)����; cKmmc}p`���v�g�&Ҥ`�T��a�Qm�����A�Aɍ����2OήAC]��}QYO��um�H�N2k;�#3�3!˨@i�k(
�Q
���6�"9�'+�z����:h�t���d.�x�YO�}7��Ԧō]q�0�٥ȞF�x��,8�mkK�@�@\0F�݇�%���<����6�H���a���;�-^�����{�p�ͯm����1�wF����!;����#�6q�N�@�&��]{jz)�ե�+u�vǫ��hE�!n��7��8��*����j��n�\��G���^�!�����(7&s Yb=�vT��?�+I�g4�{�[�s�Z��.ʩ��O�/��ؓ�!�4-z}�c ܽy��4���"ҥ�QH���+�;W�=����Yr��l�$>���Vx �l��[^!ů��f5o�������iE똟yQ
p,F�t4���8��щ�p��r
�SOjE�{O�"��i�ܭ�H,�>�A�iVCQ���o��	f�Qu�V���'�43y�ʩj��@}�,�.�_�m_0M祈�m�yZɿ&Bn�*����80�8b�� ��׾*�;"�O� ����Y!�8s���'WWL��(�H_����U��8��q�=t8@�eʃF(�� �����,�U�2 ��*g2���rSZ:Gowt���e��eh$ݼG��~t��$�E!.�F=ƈRt�;|c���>ԐA�i(|��bC.:�&��=��� �1��QE�_��Y�/�����0��ݰU�z�Än3H���G�B(�$���!�5ɯ|���~���MT@���W#z�v�����]��u�|�O	��{2��gm.y�$�OE��昷nh\Ȝ
U*���?��KM��N-��ذ�q�	�����?"-���61�9I��S��^`���bXho,;�/e�6�4[��k)ǻ{��O�_>�+)�r�=�FYʂ�.�:B�)$���6�5!�D���i�+,/5�Saq�B��Ն�VVߥ�;C��ڰ��]l'c�:р��n��HY���[�^Y��9���,�^��� ���E@yŒ�_n��@����^ޯ�|���8.�,�2�-�3tDAm.0���E`F�	�@�1�#|/�2��r �6%�%������]'�)���a�~_��?e��J��q���yH`����L,��<����M��R�a�娨���yg���:�0']��(��AN�C���*����'x�n�# �V��M)��4�80�XtI>/%o���2�@0Y����~(g��tO������>�ܤʅw
:4�;�79>��oW,�n�n��J�&{���ȃqώ���<�Q�R�w���@��hʲ���zY�?(�m᮴��
>�.pZ^KdA��<�:,��9'`�M�qS���d
��9��Ef"�'�3����e��g�-�B�vK@aC֬�����a߱�9�j`���x^#���8��x	ʭ����&��������p}r�A�״HЛ��&�$�|�����O֙������}C�0�?q�4j�n�I���|��x�U�$Y��E�#�wG	j:���D�+4����w�:
�Q8�'P�b��վS��`��})�S$촼@��N&��n���A��'3Y�}��iv�e��wŕ��Ao��ᜆ·'5�~S��M�"t
Ұ��_�]d��D"[�W�U�"�Vƨ�y�HC��x���l6�~?�	�k@���ڠ�D@�V���1�/�(�6��~����g�օrF���ٿ�(S1ng�M�fjr��=�w����\q�L(�WvB����W���Yʒ�������vWjE6���CZ�LŁiM��{�#�y��7��
~A�_Y�\S��!Vz�斨=s%��/�s-#�^`�Y�M=l�m�cčǋ/�67W��aod�f�U\���ܬ8���xW�����n�xO���,?i���h�_ ����a@u��� �Ȭ;_O�p̂Y�*_@��f-E�9$���@ w,�hb~/��Ogt�� 7�!^>�cCh8���;�����y"��>z �*n�(�M;�L�)�a�_N����A]A�J;��!�4�~���vz�5O��Ţ� ���� -����i�&����B��A`���|%
�ᤑ�JR�(��i��R�hA�َ9�'(�\��r�^+n�^�3��d�EC�E6/��w�l�ß�B{�y�x\#�;24�#���zGy���8�ӷ/W�-g��0gӼ��N�v��z(�I��=��8�a���P��.����M�+i�YAe����٥�,��'-�@\��Q&GB��)��Ypj0��ЭA�<�4��{��If���3kӌ|�	t
.�=�ޞ Z����1��(q��)���bsx�Ё��~���IKs��B䄊�i�%���� VlL��^j��7�L]U��Q�NbD�N�$�.�q�'�b 6��p��^�,��>�`P�@�H8����W��[[���%M��#'h������]��Yh��DC�#������G�	gs����ș�Bu8=��Ca�|Xx���Z���O�F����}16�ޒ�Ew��E)o��,��G%�h���kі�Oٗ���'�oU(n�\u�MCu-�� �⭆��lF����S�&�=�eՌV\�3�|��#�v=�l����	�0JY��ҀF�ϪmMY"8ZXl���:O�aH��ó�����9(K�o���H�$�j�b��v)�>q����ş���f�5����C2G��>�q��*Cpw�)���g$��4p2Ŭ�4xy�]H�e)��|yV��Ct�~^�ۈ�Qʯ�ĩE�7:蟋*�8N����2R+��9ű����.M�?ol�� ����wO9b�ّ��(>���H�&9�m��+#@W�T��RQoyS�^�2���k�"<�}���1."u`u��Gm�-��2�9*j;������ �;�g� ��Bfc��͂��}z�M�Ɏ�G��_Y'_�~Ct�3��aPϏM�k�ؘ#)�%O����~V�u�~��H�Cxj������g�.Х��cHQj��;�R�~ XFUG���P��4��m0��t�����ߓț&���z��0�� ��w�]ټ��_���6<���ǮԔ���V&9��1�-NvҎc�����ʺ���4gc��:#��w��#}/�/�B½���q��Di�mg �Ԏ�)U\�-O\M���B�L��JS؏c�VG�*����5�W2�5��VO�o�i�	L
��V�Ю�k��~0N�b�=�1aQ; Ea?�U]������� �M���Y'��9�k*zh{��#�0}L��0��;ќ��YXzxf�#g�T�$��g;Kz'� �@i�	]�f�ӯ�`S.)��ڛcϫ�E_~�g��佾˫y�,��T���eSH�uRz�O[�@ *�ॿXn�!2�3��r<�{hץ�6B�3(w>�[p�N\��w�G��Yf���O��f�&I�w/���j4m�S"�>���K��p��X�䟺�D7�z�U2�ū��m����UU�;�/�>:�-�,&Xv�G@�傔໬C\� ��~��\k�Qh(��L(�����DY[���q� ��Jn�f�V}�m|���I���Y�ռ,���~�l*��gADz3��Z�ޮK��pDn
$�x��ܯܴ5&8��u�c(H>��l�=������zt�į{Ю'Z6��lZ*�+��H�2��!�%>cn����~33)����Ç����2��^�^�͏��@�����k�	���� ����[3;�٬�Ԙf02L�ը��:2��%�ܾ�F0���v����i���F=ku��*G�����JE�Ir�]hY�!��M�L�t��d������f裂���]x~�F1�Fo�?\z,{���A��',�PS��a�d?07�Q���,��&�Ϝa
��Ȩ�D���ʧ������_��g�Ͽ�p��Z16��#��8V�&��go�:��䠐Bd���7���	\����Y�c�u���@5����"���BȚ�B:D"�8�ts?�ںG��V�YS�M�p��q����9��ǡ�?�v�	*�#��j�)<���p]��^;���g�`w�!>�n��q�R�ra����Do�QB8b�yI����\鷞�3d���d(��w�8�^��;y>{�QC�k�Z׼!uf zR��>�&���5�����r�l%>`��G\���6{>̗2}􋍱q�1^���!ԺSA��<�.5�o9��,��x��%�A,��?�ơ%�8	W��H��ū������b��q�8 j���;,+�Ӻ�~�]WiH�e>?=�R�W���*���9?;ظVP{���o:&u�=�5��6!�2���y[`�˦����O�z~��K��H�M��Q��;a���K�@�'s��>�ί�y��6���K.�zH�+b��<n)��Yg ��,y�N$�� 3F�ɜ֋�EGk�^�3�=�{Z�ː��!���X�>4����G�������ӥ�Vϸ�E~���B_�RB��$��1?�_%��U)ߏ���̇`�J6��[�v����(���4�M�re6��ߐ���6�3�&��&�V��F��/�D���"0i�U�ע�R�g�@��i��3��f,������Ll�\n�)eG�[j��B8��^m���҉"�eFx�N쒆��D����^�A��������@k7i	�wT�[bb����T��l�u�;��U��P�(�r��d�%�lpRU&�,="�<��T$㭗(Q�AR�5���ݘ]�H���g ں$ [݈yO�m��hRG��/�'������k�p�0�[�9��"f؁x��aw�k��g���<+=��>J�Ei~��UI�Q3`��s�H$[��>�[%��&��f���"�wP��[n r3y	V�y�e��r�^w � k���$��L&�`C�a)�/�`�5�ai���� k���eB��k�i%N���:��.0$gWe�M���Z���O��A.�'T Z9�a}��B���a״�3D��J������^:�p���~o#ݿ�*jH8G4�pd�;��Bf����H�� ڪy�E���-���j�j�1⇚�㿢mΈ�ر���}U�a����F�u�&�}WE�mf��Ҁ����~��f5�M�E6k�J��)�
�y���(7�gI���Bn[sM[xeLp�� DգNl�>
�a>8\�l�*'�DҮr�I�v�=��oX)��UFe�5�7>�d�c���a�<��h�v+5�l�Rf l��ġ��_�ޕ����K� g�!>�x�
d�|�1�l!���h2MT��"�#���S�´\(K7�A�b���R,�=���i̼o$z�{�X�m��y&W6� +��k�G�}�TZ�lH�_"i��ra��D����f?1���m#�<߲N����B};���q�_>�3A�v~*xj�}|�g��i~r�|ȠN�j��²�b��6�Y��P����������;�>��_�}�U4⻯w�%K߳fi6I��d�s�0���E�L�a����e��F�����G�Lv�9��.%��o���n�;C,�U�o�����l�X����	�K*��}�Ņz�2U
��}�մ������CtU͎�5��*��G�M�#U�}̺@�z��切3Yqg@Ѡre�7�f���G�'�uXlxVHYEB    c945    1240WB�W�nR��n&��(�Q2)�6��_��H4���bq1&�j&�VrQ�������)�N�-��=t�9�W/�jC�f��e ��Q�����e�)wD$�C������3y���$X����z鵏؝����C��r���.��e�8��X�>M������RG=
Ʈ��ū�o��?������p֪�Ha��r�}��q2I�h�#{5���.(�%f��CJ�0���ӛ��eN�Q0��t݀2t�{�-�%`�t�S�%�&��dr����\0W#9�[qfF��"�9�%����h�=����m�EM(|�W�����(�N"V����8�3��}��WuZY��x`xt�B�O��CV�q��B 
�.*�������>�nb�=�X>���ei���H�!�ŘN�K�kr3���1u^P�&�*�l�9�XW�.4����$YS`k,���������VT��oK	�aJ�EW5����Y�����Md��/g�b=:���i��+.�����J�M�.��}ċ�V~�S����G���N��7I�G(u`�����q��5=���]���?2�N�M˙�G�-�3>��F&���zBS��Zs�2������:C��}"yߘ��F"��w�GA�}��r|�&'��%��~�U����'Ƌ��	A_�}A	����Tjf�*:	�Y����V�y</��u�J3z�3o���b���1�KU�K�s3/ ֺ��kv.i�TI
�{����ՠKuj���Pyf��d��N$�:/�_7rV٩D��6�<��{	֣�G[߷d��{1zR��(H2X;5��E�|�{�wlAn$'�󸡩��}~��w����k�e��,͢�~ͨ��������5���A>���#�ˑ�}-݂�:��}�[i�Q��$���We�1��ug��1EZy|�0��>�Q�"jo�j�9���q��b�8���K���$&���Fs獰�a�"�x�l)'�l���j+�Ҩ��d �WG�8��q`)m:��wg�Gz[���\
����Y����!�!���:���ho$|�ôIj~		��8@����{hߌ~��aH���C��{Emg �0biΔ{�Mz�����",G�8����˚
��|��fx ��]"�X8��y���;�.0�c�S�v��n�>,����2� '�����IQ�^dP�' �8�0`^?
K� Ŋ^�h�� z�uw�.�?h�dt�`~3�˾�ڈ�2��}��Ò�]{_��5�	ו'����\%�0�>Ԧ�Q�v��Z�糪D��2(�]ٗH=�Q
/s��6]1�1./g�"�G��)�6O
%=:S��څx�-~��s�»!H=��|�};���*]����*����ݢ%m���㾋�k���#�72�>���d�� ��-�L�JI�݊ro��1IsU�Mѕ�
F�\O�3�D!�(3�D.O�kj��5��SQ����SR�Uy��1��N��"�^�DD����\ B��̏�
�1�>K_<{fπ�-j����Q5�{�KJ�_��1Y�^����6����N1Sb	?��\�]�p�ϸ�?��,%����tP���j���!PM�)G��0����b&*�ӈ[���SAS1d�`#��Y�!\o�S`�ŢL�r�"PeD��v�d���r�8f�D	k����I�
(\3���>I�Ԁ6��ȩ��uS?�ߐL.-tk��2�+�9����^7�62�~�hT�Z��@�4�-����~��v�����3��p��[i)��x�
�'VX��+*�HV�A�.W|f
�����JT�_򋋸��f�c
��C�OoYϘ���axy�_�;�4��X���e�S����|o{z���I�M�`O#�V�Δ�C���}'������lk���!���M�7���Z
mJ��b�n C����N�����-~�̾5c@G�O-�S}' ��D�� �ɰ1��Q#�z�8>�"�p��`Uu���ڰ[biV�e9N{�+ߟ�D� ��]����=���}����Ik�M%�g5����|�;o�9v�xtc�H6_e
�����٭9��M�2��u��GKs_�y'�?k�)�,e�u��f2�|(Жa���Γ ��I���ƥ�U}�Я��_E���J�"^b� ��[�5Y�L�Tؘ|퍶Ս��P��7�����ۈ�y""�M�7��<����?�b;b�|���2����K�ᝯ8���)wr*|��O����T#?A@Syj�������+ޓ��$C�i}m�&�R�,i#=Ij���"q�ͬ�P�ϊ��x��z�cV W蜕O�*��<���M��'�x��o=�ܱ%��;ʺԟw�Zd���q�I��_!���X�奊��3a�R�٬>��	�	�Bn�=�M��3�Dv��Uj�՜p��S~����"�{K(l��s�>D�G)ΆrhYN�u:
ެ�C�Q|�4'{��¦1̪� 1�D��n^�t��C��- ���r�0��B���ٴMR5�7�v$��0��T������u!]q+;E ���V��K).jԷ�뮄�k.�1:zk�І��K.gf�w�M���S~)i�D��O�����'A�#�o桙�10![1Zr��v���c;��p=��(ۥz��A���[&/<,�K�N��߽l�I�}_wȡ)`7���g��uPt�=��#x
����د�|�0�@f���EQ�Y�0���[�?��ę��󌖴Lg
F́	���hPn�=��,���\����_�8ֿ7��6�|�5�K4��k�?Y֯EBE�#�0e@�d�<k��a��.��M�<����s0�X51v�[d�/0TL�����8�mg�9��t�;ѝ�vGQ`�PR
^d���@�Ѧ�Va���I�Ӻ�t�O��/"d�o����Vw]l瘲f(�Zpx��Zع�m8A�y6�6h�Tz�Q�*�r�����\������OZu��=\[��2�[�wX#N��3(t;W�z�G�2&����OK.&#��b�z��3i�����+����FC����3.Y֚a��-ɪk���
�-z?�/�G��?1,��c[`�ֺ���M|cO�KXquTұqD��/2<��\��k�Iޣm����L4�&�5�� n�2FZ7�\�q�t���̣��j�H��'��@���I����<J�=*��`�N0͇F@��Hu���9Bp.k]���T����5Io=�:��L�>��ܱF��s���=	Dj�>��D3�{lsw���������֝��m����	�j�M�ߐ�X�������l���u�z�J��u|6AJ�p��S�g�� �j(�Z���y]���r��`�2E�&�Ƃ�V8����n�k�S?�)�/��ؠ�s��N��ly�ie�eAQ��f�tH�=�[���6���?�<�E �vZ�)�j�`�G�u���8�MЊ�n_�iR�����<{��f)���d�f�����.��R^\��ץXO�O�$�{��L�n�㌒�M���T���W/j��9l
��O{�aV.DZm���l�h6+3X�Ƀ5p��~R������̈́v @��1}��m��ϟ�v�;u"�g#�]US���1[Z�?�M�*	u�O!��l}�Qz�%�ҜjH_���%���+߮Dh�@/���,�E."��>������o��U���[3f�M��_k,��<�E?9�޽w�)�m�@$���7�G3��2��c�>�pE9h��Q�1�Yu�����*�I�f��&y;eܿgy=��Z��A�T�4c�h������b�8�x��Q����b�<�nu��Z:BŠ�
�ElL9n��/SE�MV�3�I#~h��4�	����v�L�<&������R�uCLw����%@|��ׁ�Sr�����ZK
L=Ç�9���?"��(�=��N���x���,��θ�y�4M�<��;f)f�ʤ,?'h�]�ӂR�O��{�"x��Iŋ��uK�E�Ӳ$�H�_3�:������l�L%�"$ce#�@�����ʣ���p:��A�N.�KdC�"*+�yu%�-"�]	KE��!!i^����n �	�&��#4�l���7�(�P���z&�-�#�s�EpST^���u�o�Cw���Ïcf�*�2�_ۙO$h��y!KE���R�Ȏ��`�b���s�K���+U0g�'w�Ci�M�ԌU�㶗��n�o��ɲ�`C���̺z�3>:J����c����N�`��;
z9-�":�i��Q���IP���T �vv,&���='зoiYĶ&�y�ɜ�抮�l�w��L-�D�\���E�����c�β�_�`���;�O�.�ę�@�	�G���%vy��#}è[ ��Ӭ�������a}�� vK�
���/��8*�>�9�7�u�;��>!@#Ӣ�,�%d|�
�b�4�=u��y|.��T�g�w%bu$I�*�VɝO>;^��Q(�07b�q��"(5��r��K��=/�		����������Z�=�9ʞ;�d���B��a���(��{�����n�x�)1v��"��]�U؅+ڜsO:�2�L/�&��u���a���A3��s稙��ց��9������(+��H��&$V�y:�9;M�i�8/vh