XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��B��-�v;�]81��j*����8�yp��+�i�:	�a\`�A_&����_�F���]'����V���_)P<N��V�;m0Ό�NI���VH������߂��`m���ܱǌ����A�(]8��\�b��7s�*��*���]���0Vڠ�3��t�/�-�]x*�$.W6�4�>�V[��4n��n����pH�6.�?��H�ڬ����)SJ�ZW�M�
��{k�E�W�O������vWoR�Y)o?�6�����m���`2�J���2���'�f���aoQ�����j���R�R�w%4)���:h���<#¬�}�+�<G���j^Ӷ�jaᔦ��Iͭl���Ʀ��SC����}�_�/���;�ÀU�Hg��-��;�|��K��*���vF�d*�(﷏�|�T�|�$��屪�>LB6S��p��Jk��� 4<��G��!�2x�1\�ػX��}X�n�>g�l��D ռDe ���m\o5�I?��-c�����z'���l��4S��ʱ�t�����"�=�[�1+P�˛&�.�K%�X�:kE����6�c �������D��X���Y,�#�-�?D
B8z�����9���Ƨ�ꃭ�%����~����f�3���T&N̚�������'gӁ���~��%�u�f�e��%�4����xܺ`*��o��ɠ"�\�����\��1 :���M����"�rBi}��*�����r�1�{z�N��+XlxVHYEB    fa00    28d0kN{^�^����מ+�J���g��g�w�c
(��
�"@V���ֳd�3y��iໂwO���$�<�Ov.<�>얪F��\����B4[:VMq�K� ro�6�L�9N�\��I,fk���q�<��A#�Ӫ�L�n�U��_R�ZQ��'��ډ��0��P�!�/9]]<��#5{܊���� ����GZ0��[�p�pRao�Lx���\*���J�S3����	����5"��":�����xj<t��uq�4���멁�Ĺ(�X�:<�KR/?]�nD��i}RO��jQ��#��q��|*=ȳ��#߁f�v%F �M������{<�N��H��F��z�)�����&3��T'#Ro$hg��������OՋ[�����;�>�^�����o�΃�n��qb7/H���\�
4A�UC�2guo@�4{Ȫ�"��|��t}�)�Pn/8]ɾwP�*�؏nG7; ��{���S�^�qAZOrl^�V���6x�W҇hSa>�iVYv�{q#!�F��Ek�C�<9���J	�����H�An\�4�hP�6T#�1���4L>�M ��l����,�3e��=ѻp�1!�9�;!|��;3��7u�����#ĉQX��7�����'�#d�����#���ߤm�F@&��=Z�XI4{� 7�h�8��I˶��+bE^�=n�����T}:+� �b�2�ka��}������`n��:�qZ���.l�'�8U����6�t.V,F��'�;('8OBy���+�W�*J�%�D�nH��sճ{f���W۞�����P�Y�!�PF�M�V��4�@��p	d��FT��l�Mc<�
�N�T03��*"�e���������AZm_\I�9&�`��}�÷
��('mʻ}��j8Z��ck�nɆu�����{?~C�MԳyz@�'O��.�^'Z~�c$='��f���JH1.j�|�G��Q@d`�uC>�Y2Ɛo%�D���#��,���&]J፾c�����.=�م��Y{���\��8% Qk�b� �.��-��˫�N>��+����Q�̒�}ev'��)��`˕+4����4���5���2��Щ�E����F��>V91�m������b�BP�5�WYu��v��{�r����Z�=��^	B��1W|2�o�i��d�2b�ʷ�����[�����HRd�6B�T0gq�_�vDu���ݔ����tk��}�Q�hC�%3w �d�'g7�k#���.c����z��<|j%v��K�$hrV�ڛ	�����g������RALѥQJ<}�4	h�AX�pLc�9���\�t���ƨ�;�u����{�u0v�7rɻ(>
�1��κDB�9%����~/r�JI����׍�_���ŀ���!��i�y~C%��[�dC�UA�(ڞ�B����zg���,�w�&&�E-0��c��U�cr��B$�I�Aצ�46�
3#PQ㾩�H�@��*���`ڒ��M5$5�e G�h:�����wh��Fn��DxR�vW��<PN���w�L ���#)ĥkgEpFp�lf��<@ ��d����	8?�m��N��,���_��i�\/��w~/N�i��O,�d�8�Wu٪����y,�}S��&բɻ���+�� N�[�҃��o-�cP���\?4��;jǜlÀOd R����O����A$���ܟ�+��`%��l������\�C!�ʶU�De�QMS[5\�#��a6��.=��?�jю��wĩ�
���F�.ӿ׵P4�S+v�}X��_�4��a�We&Dƥ���f�i�ʿ9�w����hA�'���ŗ��it��S��;�������|TΡW�R�7JZ��\��&�"e�'Z�)�c��;B���~h�'��"a��@W�-x^�r�7�N����sdw��Y�i$�kh߁"v�)��Y�"N&�7��:����B��P��|@���|:�'Tr���?�w��ke�X���&&�MP�{��&��;�0����g�<9!m6$A}T*���U��Z�
�����
�h�5�2�ʘ'�"�����]��x���.g:I|��`��B{|�4�ȣ�,�IU~�>�¢�G����(�o��~�9��Z:�]�楂�S)e#5����LJД���"���UW�ɺ��!��ş�W�,���*Ņ�d��e�]���*��Q��%��w��p��4�ҎA���,����L��_��H<�Q-��S�8Se����I��o;�j!�������=v<He�Ab�"��2�`�v��U]���.��}6ý�Yc�r)	Ō�䂵Z��p�9�5*�@#pim�����x=�EZOY�u*��9K��t�k�����9M[	�e�,B��$�3G*����,���@����C��Q��=�u�V�
q��$-�c��UٯQG;�1��V��S ��2��rn���ʃ��(���B���T�[ƧHbF����g�r�q���ۍ���Z[�͔�̟]�Opy�P��x���xA��M�C?t�o�˩���|ݜ����Bh�Dٸ<}��)^-Y���h��GqwB�d�5K����8�{�����Wo�*"��2�!2�̉����p���+`�]�#���9?'���k�O�-"m5���&>���#'�1[�?�H�u��u�DXßF�
��3D�n�u�?�x���ơ%z�_�p�{b0ު��,y�y_�L�8T�)����0�[?6p�G���m����GX˾C���PRejEA��2������m�k�;�7�DF�?h��g4�FSDQ"�b�=FŇ��IG$f���FwM.f�2m��n�����ҡ�[����}ٚ���:=z��˝d����/�1�y����ѐ`t�_غ���1ϲ���䖑����������8�f������f���M��
�ړ���r;����&}Q,��W�fhC���־� %�9�O��H+Kl\�Y#�STo��+�l~�IN�0����z^�
-i�-n��W��y=�_1`_��̜u�/�u-�v�4[�YL��p���bw��7�J^*��xꣾA��>�������p�k�,��	a%�DSvʦ�Th����872����E�$��]�R��T<�SG�n+ڀ@��
g%R���ƃ�����-5�eS)ʎK�}�z�]�����!�iQo�z"�t�� [����`�ő�U��'���1 �K����=���8�N��A�@�7Ѷo��
wU�!_�ŗS.��� �>���Jp���	�����������T��_2m9[+�<�I%t�Z��]�r�jQ�d[3V�(��fY%��yV���{ۤ״�q�R6&K�ke������� �v��T��
Ս��_�*����!=!�z�]���׀�'�e`xpjÚ� �Q�6)-%?.Sc��t���=�<j�����k`��]���t�}��]d;@Z#���@��m�mNDɽ�i�3�OT~Ά_yb0�+�2|cߚ������D������a-�<Q���+�nP��-k��܌c� �,�_'���Pz)�������/ݮ7$�E�X�Ԇ(��@�wg5�`�q�9���T����ܺ�\��u1�T��<i����D܇���]?��뫨���o�pa��K���zX�����"_�����QZ��H�]|7FpŢ+�>"L,@K���(K�Ɗ���
f<�YR�QPJ3X�h�9��\�Q=��=c 	�J�����DxAZ��g���&]��&D�T�X	�D5̠��Y�:���>���̤�����'%�q�S(�� �1E����'�"���AI����5
��!�}Z\���0�Ce!m�q������L�,����N�����-��ӱ=��EH�&����ke� ��<9J�S>�j��6�:Y�������V������p�u���M���5�粆C�oq^����X��^z)x���hK������a��}n	~�$"��yu1�=�����SS��C���z�'OLG���,z�T�;�|��##�c��!
D��23�y�3J�K�M��-c(_��}�+X�/g�ي,���ϡ��B��귋�/��}�H]���p�E>@.��ˤ��}J�� �.��ݜ/���4ג��E�Y��x-�DA�<�Ԍ�r�;�7+�E�D9�k�|z�7>u�f?�f��ۤ�Bu��d��>S}���}�� ��?�;�~#��/�����:�N�mM�������֟��� \Ig��$�a��M^�24gO4(�^���Y��/\��y�Goҙ� �r[ş+h�#�m*C��
I��;��!: ΜE�xQ9!H꩑{s;��|wd��K(�ٱ�j���nx1�i�t�T�Fd �h�2�g�]R�_�Ûkxu{�3�j�@����(�M&��w�=���D�C���9ٝNC�m�s��x���~ɚ��YK���ug�$��A�W��}��?�a���U�d��H���4��p��阿��Q���=��;���%���qN�2D�B�J��w�}��P?��
�i�m��לW��N�ܶȳMo|���va�I�hq���G!�al��=����0]#�����ح�H�U�R>�̍J��9�h�{w�T�PÇ��$@��	r]����n{�]��6�Gް�����?�qZR�x�NF�k�gS�<}毤��;n���l�A�4o�;{Ĥ��@���'��X�����#��>��8�B>c��E[�rMY��(��3J�]�.L�Ҝ#ۻK:S��u:i7l����%��}�ui �2�s�z�M�w�ګ����Xv�L(]��aZث1�X��Hn��EԣZ�͉h�r�'�9�]��re� ��M R6���i1�y�UJC
�����?b�� Y�]�(�YD�De����ٸ��^�z�U�=��4P�^��d�RvS�b�E��T��-�R��k{�.K�d��9NE���q�VV펰��X��+f�Nܻ]�Xk�����39fʄ�	�'ړ�5d����srW<K5K�UJv�����IP�>���X��N���j+���YU{S7�)��9:�-�-S;Nї��x���i��v*ߞ����o������C;V=�;���̾�f�
/UJ����^���@�yC�1�v_�ƃ��m�>)����>J5+$T�K ����`�]a��BA+'��8�3�j�Q�K����3�X��[��6�,��'`�����4a8����r4����!I#�ҡa��+[��)?k���F�8Q�t��yO�n	|j�Ŋ
O,	��g�i3�W-�����[�(ፂ��@^ov8�B|���Y���5��6Ƅ	�Mk��1�5����BR���gE��ʣ���nc;g�Ϛ�ʱ���U$�wAT�O��IE-!Q��s�`h0zRAx]j�ϡH�AvGEf8W����G$E�ߟ���]���LC�0�T�S��d>i'_j�FE��*���ħg�
PB�u=�����=w�p;���/����j�����m��Av�xwP�glOSu��򄄀�p�_�`��gz���P���_z�i��;�y��r�;h���QwШ.�"��G�z\F}d�JJ�P��G�����E��Lj\#���*6R�AV�H��T�� X�Ha��u�7�n��_���ye�>�-p%�H�������CMzr�D�w����kr� %��c���ꯅ����3��˹ڢupn�By1��P!���⥯��n���Z��Ke��Ijb��Y�c|�����3�Â���*Bze�-�R�G9i�
�"/d��Ɓ���d6�oD�{�s�h����<GC����J؇>��5�/(ԅ��I���1��n~�3���CmБ���.��I�Qa�Bs���0J{h'?�v����H����l���l��x�)�󱵡�����}<�Y�M�bp�s�z�N@Uf�G�?A7~�=6��Q�� AAHwOD�^ސ
azc�l`C���Eh*ۤI�>����4�[8u��`X����]|Sx]����nO��X�0�5І����
|�N��г+]v�dԬ���W���o�%�B���:���G��g(�>T,~�*p1����8*l�7_�S�h�S��O�(����A�W��c�S�JJS���=$��c��j8G��c�Y��=.׶M�>4�6/Ѹ���>��&��Yo^x�k��C�Ӟ�"��jS�`��sf��}�j�ModaC����6:������e������,g�C@�r�(z�r����5O�s
�3�ÿ��IA� ''�!)��%���)nr��Rȕ�2��r����m��5�4h���C�س
��`�1�4���Ko����L����� �Y�U4(�"�E�#��q��(B��(7�$/�~�%�
J�����x�����O��.k�\Ѫ�0(�V��YV�;Ѕ��9�?3 / �f�b�^�l_��b�e�o���V"{�`t8�.��D5��f���m�IQP�Y��S�_�Yy,���n���Ƌ��Pqh�@io<b�1�.H�Mf��E7(y0���#��X4�����7�d{��I�tc����	�Y�G����#_�1�_ BfDMI���*��B�e����8����$�fqA�P�v9��[��r�=,��_��Dl:Σ��]���v���ԙo��i��N'����^����Ŝ� ��_��E傐��2�)�s%+���F�z2�U�	�˕��ȃ�0�m/��e����(4��P��)�ո)��p2�]@̳�@T�c�m�׆����ΉP��?*�찂M�����Ń\E��#�����7������
T%�>Y����4�v�Dq���;T�#v��x��/�X�F����{�/�a��G�dR����'��t�=�m���b��x��^6I��U�@%��9�]��%r0K�+bI�q����d������^������G�����eN_�p�y��F8���;���Ұ�0�!�Z(��y��y��Y���.)6� b��Ds�੾=��}����!��.y�m�qu
�Tb�b�H�~�F[0����ʤ���y�]POA`�EhL�+E�Fњ��7�� �Yg�*�'S�7����X���B�Vb8�����S�~�	pJ�����ޓ_�R��<a� ��袒�l��@R�I�`�L��,[�522�w@w-/G8׃c���?*_����������j�g3-���(<�͕_/S2^[B�C��R �?�W��4oL݁�U�f?B�̍d���b�.$6��C}�i5�:�]�L�$���/;�n�?����+,�t����@8�_�� 䳅����̉~U��̀����	]E��l_Y�h��i6{��I�'g}S�dZ�.D�X��e/�ƹ�*IKj*�O��ޣ�����r�֩vO�`��I�@(�Ï@������p��s�Ԫ�ʤ�4�J3�������`KC�Z]��}��y��};��)��E�N2z^��N�Ǻͯ����_�=���Ų�� �?�є}�ڱ�d-KDQuS���2��g�N�d�Uv�If���]\]�sumG�N�������W����`��'�+���4�5e�r�_�ES����Ĭ�e��g\�a&��1⋩��D�e�(�fA����^��?�\CƔl� ��|���S��e[D�#ap "��m�9��{lo�5˜���̐��	A�:$)��,v�GwL�Q��Ē��4����{ep�.����RϘ˭��,��O�Ȟ%��9 ���}�aw�e�q���H���P�O#�[:$~��G�c��?G��~ �e[/��;~���T�\Lݺ��@��UԻ����M����Q9�B=�g�~�1���^�C���^���?v6�D'yY§��ި �k��b�z�/ ��O�V	��5��S-��0���P+��0��Z�?�����e�X�za�	Ө�<��
�i�c�Z����j��v����Z�}�������Yٓ����b���5����Y2鼒7�K�fh�@�=*������,'��]��υ�n�dd^�Q�0��v
T!���G���j[T���z@�z;vˠK��f����c҈�90<�@z9���9�j�3�u�C���"�!)�K�(7�i��)�\1���o 5�ư�>X��>BX EYf���-G|�ch0u�����%ieo� �48�|���2h��+�*'�����>���5�g#?:~3��\��N�g��K�ʂK�q�_��7E4�W�b&Eb�	>���zt��Ò�Z���Q덟�"�ꇩ�y+�NP�r���^�sn��X� �:H�U/H<�Ꜩo�����B��3+a����A��N��o���
��rR�wzW�D�$Xn�w/Ƚ���>�H5R� �(�-h����y��qҚJ����D�l/��	�s.a�2����B��D�xe��/#O�J����)��!;�C�+�� �(�ɡ�@�NH���r������c�:m��y˭Р�:v*P�����Q~ �d~���qV����Y�D4Jd��[���6v�?5��LLeN��^H�z��T؆Z �׫pqW_���L�K���hk�L�}�C^6p;��}�`�І���c�'%�L���'��m�F�x[�	�%_����c��2kJ�H�P�[|�{�z���
�ٓ7��!�H>ك	E��gb�>��h7��2�w����p��R�����q���uѤ�����5�6�2@,�M�08)�x��hq>9*oBJ	���)�/�[��#g���H=�;n9{z�НC<��
K3C>�x�׶�ԨA*�R>�;����h��������c���x�9����h.��"�.�N�e/:*�~<z�8<Y#�`F~���ýIY��S�L_�<�!ҌZow�O�2���N��tj�qP""/(�a�O���*�d�#�/h���F%�ý�=x��xK�񌃋���-��n[[�򓧁9����m����韩 ́�/@ʈ\s�m;�Z�Ǔ@N�ñ�
DG(���Z��5I�r/L.����4�x���7��8�
��>�J�͞Z��oL��eGʈ$TI���e8BP�k��Le� �Ѥ�@��?J�b�d3v��\i=	.[h��Z
�x'[�e�ƳI$`���|���uO͚�i�J01�����@���G���Y�L� �zu�/���T�8j���_�P5$p9�Me�? �}X.!c�/�g�<e���Ϛ��>ߒY�;C=��e >�w�f�L�{��!->�dK�B�{$�7
��ڽ��"��d�O�**P���OVu*z����l`'Jô�;m��Yy}X�������x��k�U�
��5�W`�Sm����p�'�&�]��K��G�0X�}f��A�#�_6{�8���e�~�$I������U���5c����hsA1ӂj�B�w�H�A�C#ޫ�7���M�¾��ߧ��rH�Ҭ�N'pP���ب[�urp/���y+�d�p�̼	9I��%E9Qֽb�:Ŵ���}����	T���ť��V��;;<���6�.�c���t`��Q�#�;8g���J�mz��֡�(f���K�1^��h;����A��y�Z�,fy�:8(���G��7� ��5�c��MF������5`ŀ`DRi1x�kQ�9����(0G ���,��_'��$;K�+�w����K�`V�0��d�7��,o�xN>�o�{�}�*��@���)�B��c^2����{��HH��L�yRM�^��b5���_@k�K� T�=���}=4!o�^_���?-zbAJ����6�U��+��1UZ���+5T��)D�:&Ϊ�*���}��b��n&;Uݭ��8X����wWP��8� A�?��W�]�L���`G�&���דMdGH�e�fy�����U�ޗڽd\��(D)|yL��Α��,�S��|I����0��:
ic�����'�_�p�9�������#[`� _JK�L�/W=G�4��������يtMp����w�@��E�r��J���u�T��,ƫWV@#B.�7�<�^���,�FW;qh��%�{��Pƌ���	�������s�\�0�������QI\��~�K��~�3U&v�N%?C��v�M^
J����3�=:�;���<zP�{AY2%�uud��_<C>-?�
$<��
XlxVHYEB    76e3    15a0�j�9O�I�$ʴ���1RL[S�R/R.�jT�so�'&xΣKɣ|hu-p�뺳�3C�hc��b�[DC/�c{�[��!q����Y_��xX`V���l����A�(a0l�BWg�+|���S����P`��W��I�&ۗ-6Kp�B�,�	�Z�j�Θ��1�������p�G*�AW`z�/>��!���y"�>_�R+
B�T��>M� ���y@!��I��2����/=��D��[����]b��@����Ψ����i(	��T�b+��F� �bH�NfT
Hh�[��/r����L��$�����Y� h_�Z��F�K��^����KR�������b�X�Y
y���8��t�_x�����M�9�\�>-5��i��E��L��TKԤj�fL�����W�o�I=���EcKd��cyS��8J	@�W)��u0y�ϒ6����bs8�J�<ўU�Ŭ�`�	�������`�'*m"��zH���'~>�m��@�'������XOA���'���a�#RN�k����(�8Ǯ�(�:�kO3�sf��]�;��lhj��(���O
�<@ �'��c~��0 �&�I��爫�� �[$��u#���1�]i����,��n�D�И��p����k���2��w����H�Jk�=���ܝ�GE�^�NA,��Bܒ��}(62`��D �G��WWL���eC��(V�|��O��P��в��Tmy� �љ����%*�`zX�ᬅ�K!�HS�����Z��[8�˳:CQk�+��i�&jO+-���'��/C�aFzGLÍ>��7��������6kx�X��ߝV��s�_�A�~�����$���$�A2��'V���[����w�z�4?��82�%k�Nd�a��)Hr$y.&@����S�����~��r���(M	������B�9�J�И�젞C���QZP�	0�Iȇp� e�vۀn<g��,�=sg<wǒO��e$a�X�~��c�]bo�:�n��.̂k�����A{|,����i���0Ca"���1�rX�R���t�i��vM�Q[��9�`�^_S�<}ΩS��(��2>�3��>��������YI��C��&<��R_&��@�P}��|��8*BF�N��	V��N�Ny�R�&N��g���?��{b�ᣂ�)	^-�v+�TfԬ��c��a�i����C��F��--�Ý�ZH����z���Z,+$WI��F�*��MN)��*onI�蕏۶�I��?|@�I;����5��J~n�N�7D�#<�zO9\���a�VnYS�Z���T���U@��9�،}ut�[d6��c1�۬EF���_�2[�x�y�ǒ���^�"��[GۚQ	�k�y��]�����������|L�#^���ξM�J��V�-z4�[	�m��;m���f��u�Ŕ�=�z���9�3~,�8MHՌ���G6����0v����s������P�f+1���n�c���/�NX��g�\��E��[<��m��6=�d�t�hU��g�j�t�3��F
̥ ��-�^���aQ2��e��)��/TP�������S3�5��j��0鯤����K�.i8�~���1�1����j�+�����%�Ç�m���_8�+�qM2ڭ[��懭z�[BO���ǯ%��bg�M1[:x&���k���~�8-钬 �Kb�o�#/�R}I�zV��Mo�s���|-E�����#�"�����_���戚�_�%�H�qwB7�a+^٧M�Ekr�ɢ����2_��:�]�N�$�������@'�Tk AH���e���"@�3�4���.����@��{���RPV�$�� V��0g�.37�`[�D�.T�`��
Ļ������U�1v�X����:�g�v��o�l���I ��KQW�װ�nn"v+w&��-�(��a��7�� ��M�\�x��1ql�-�k�Q$2�^Bf$��Q$g1��A|��%h\"Γ����k�l.�B�"�-��"w�.��Q��@����9���)�2[�_�U�#l L�,ڰ�U*]ɱ��3��rD�z���/��G��U��S�����|�O�׹����"h�e{���0h��ݱ�B�����#��}7@ܥ���N�Z��|�9�Pz��!2���jj�y�����7�7�Vl�Q�Dا��ա�!d��F͘�,4���,g���6I�{�E�t��}�Vn�?�	��bC��/���A�3s]/6qɳr.�pV�+��I����T�|�	Le�S��u�5����w����^x�	C��nk���7veܑ��Z���[y&�Պ�5�EjX��u���Ei�n�L�iв�a�N��Ѓ�������1!�t��#��4�$
��ŸSR�Ls�X6�.�Ϲ֬V-=�b:h��;Mi�{W��L�[ﻆ�9�0pE�Ұ\�'ؿ$˲k}c'��RR��F�E�pR�|�uXn�龜
O[��i�+�մ� �ƭ�Z�P��c�����&�^��i��1$8��8b��>=�M+*�C���<a�ȷ�U�V<u-f��{�P�Nuz/R�a��O;:�?a�-��`v)�w0ё!R�Tp�����C����l`��R|_ZT�?l��$�gm�E���vO���6������9������LUw����},��A����C!;�й�1Χ�XQ�b	hMD�+ ��rC�xG�E�2��w��g��A��/Evr�:6�N8�T���u�6U��X�����q3�㫻h�������-�?�M7�� B��Zi�x����Af9�����H��+�óbE[���{���	��6�;�_%��7���]�iKJ�$Ӻ�̀M|��$�U��B�Q��·�5;|��s>kzщzE����n�|.�!z��'>&�����[�ŭ��Aj���uD,�28�r�K����X��9/<��j�}`p�h.�⻙�b�%��ʜ'RM��g�fRȁi�Y���SG���d@ptZO7m�S(�a���;��#D���s*����Q�fo����d'�,t��1�����M8좁\�!��'�v���A��P�������u�~T�� �?BFF24�J^K���";B���MWnH��fu��CDw���Ic�D���Dhz�At�z�Si��0�ۛ��]z�/Y��\xL�nwԪ������r!����zY(�1�_	l2 c:�9�+E�U����#^~�_>���]	��k�ߧ���Hƾk����E�5�$��?�}�3�M�ٕ1���������Q��1�GÌ�yoL�����g���E��p>2`��#�m�繒�&�ި���M!���
g�^� �<R`"IW��~��]�3�~����L_!}i(��*|�>�Z�W���.��%Y!Ú��@��3���%�������V2�K��\�ȠYЉ?髖�=��n��� ������������H<�������}�	�[\�&����:��[��]ZY�
 wo
�լc�TvlAd���m�u8�ۺc7�,���/��<\dpj�+쨟k�{m4|D3�r^|�
M��b�6�Ϻ�U
nt=�;�s���yX��7�:ZD�@���.��WD9�%���@)�����pr�S���ޓM}�WŅhu���[�?�����w��Z�j��9P��nG�TCE׫��ֽ5@}}�3I�W};� �4, b3�zK��$�Gs�~�D�d���3��@ӛ4���N�<������b��eQ0	�,7�)��}����/$������]~7�+rsr@�C���Ț��@[ �x�y�VXm�U��s�������4[�tˀrZ���;��]����2\j�mwVp�y�
t��-^�Y�"��ƌ��5Z�<�v�1�6rm��:ay�s������@q�������k&i&a��~��8y�d�Gl�|ڋϘ�!D�pR���LP]�ޙL�)7�W;���$�Y����b�,1sc>,|�1O�D�l�`G��0�_�+��[�ϊg��~"���7�K���w�5�� �� H��8�]&�Y��f%�Y-�����S@ԾP:UkO�]����~����9Qm���Q��s'���th�tdj*�;Q_�!о���4�!~����r�)�����ow[Ҡ�����J�# ���54�'��YQyh���;_�;��e`�g(���w��X�,W� <���}T��d뾡w�L�t��|�Q+�3��r��g�eȦ�Q�ά�"���P��v�bY%L�ߎⅠwi��_���2E̘�F���� �&����i}�	q��c��� �5���%����*�># ���.ZZ��j��-�➾14a$"���`�}m��Y�?���ή����M�l��^q;��}W����O���& �!_�{��r}�v��Jd���[�&��	��6�<�p�w�0>��l�NO��4��F��4bT/��R�g�\��e=�%�_.��>(�i�u��;��6ϼCa�q�1ܶVsX�:,ZO���;械@�\��DH�Ż�B�xg&V�f_�9�MA�@�W g��]�,*Z��7A��ǱU˰u$Nv�3�sA
A�{)�"s�4ԯ[9쇃�T-��I�)&ͪ��IH)�.����N�����EP������
�� >>�zh�0����+v�0����8��%���h��o�f��u�SF3$�1�%�p��^G�x���N��ۃp���P�!�uk�-�Q���s3�c(B:ΰ�����x��|B�يM>nԩLW{��IGD2z��8����#��p�3r����t�F����[���y���#	 ��+�LM*5[Jw�!
�A7WS�ӛ�|}�����y��M~l�1>F��l�OJ�Z�Z�� Ǣ��KSZ��)�>=OV�s����V!�kè��m*c�X�����uks"��x��P��f���
��w�V���q>��[DD:���or�-�(�4'�k�$���ѯ+�h��O��n����Н_ GU ��nٮ`�����f�8��;p`!����jj��i��- ������
��\�����#�bDǔrf�:�}J=�O�t��-Qd�I�o"�F�7����sNdy� S�����&��uI�&� ����`���MHeZN��2�L��:yE��D���=8�%J��H6i�6���/��w�V�7���{����Hѯr[�؋�|H1���a�pōQ�����y�������3��ܓ��2{+stW�vs�}�\� F�t,�r���P�h�x8���3
����%������v	k@q`���˒x���3О�P�_?߃�$��X�툧D}/��y�~As���Kޚ�~���@�?ل��3