XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� .eEt��SU����.7����. �,��&D=��'��깱mg���(q��g��
�pt�@�����s��F���J:ӑ]O@:����W�����mbԫ�bL��z�jCI2R�̛����-�^����m(fUo��	d{�Ip�L*G�k�t����]$6��508��Z��>��r�(��w�./��v֯i��>'��A ;�Z��/#����g=k��K	󲬹�noN�U����l�0�ӏ#��G]���
��E�^����G�-4�B�%�v;q�k� �-EUwEi����*�L>��R�����Vu�Ņ�{P�.̆���������Z��߆t�q�)e`��l��Wq�����*;W�����[�*G����bG{G�b˂T��PI�ADi���Ý`��q��˫�+�˹������: H9Y��$ [}�!y�4�t����do\��Kp���2�͏��1��@Y��Il� ^cS�4�?0��U~��)H1�}Dߌ9�P�Q���:M���Vލwۍ�\v�ӫ�Ʉ��{��H,De�T��;Թ��D�\s�S=xl�Ǔ�cx*Ғ�����5����U;\�<��W�c`�	�;�^���p�S�:�^
��Cֆ�ay2p꣝4W���z��72�
�(�����ŗ���-hy�@3%kR�֏:LJ���Y^mt����q����N�O��}i�}�;�3�t��:�x}�#�1~�ktSE��4"W��F����xOϡ�XlxVHYEB    117a     710�kH�R�+��'c�d&�lGJ��>7g�"��+3?����
�P`{f�ly?%�^�w��fvn�V�5xۙ�m��=���ׂ�!���Ъ�y�n�]�<Z�}Ni��`N�Ŵ��t�@D���3�ڈ ��e��J��~\�ϩ�=�6�^��&C�x�FjMf(T�8T�G�����I�!A
��yЧ�I��c�kq���5b���ƍ���/�;,�,I���}���^�I(�5��yD�/.�P��䯻f�3يr\�[�����#��9�z*n7=�L	��"er�a{�m�z?E��8
�GC���Q���Vp������O�I���Mv��@=.Z�G%,0`�_���Y)L�]�"�K_�뱱W��ԈDn�c��,�1I�8��������a�X��ٸi�U�kw0L�SѬ�W��b��A�i�+�=1�jL
�R��U�|��Q�k7l`��5clϥ���Bwb۲�L�ˁO>U�Z����E5 i2ۍD�k��k��	@n%�8��{��­M�D�5cT'�&|i�꾆���_U]m1t:F�ͪG�V���i�&��Z����K�F3��^���@'�(=�K��D	'z�F/9�)��x�[�ȅ���|4���(�f��r$�-���YBx�W�4�נ�N'j����f#���3�H[��F|Ml`�YZG�7#k��^����җ7L�ہ�ܷ5	�}Wm���oCF���j!F;l{�p�Ѩ��Ε���a�,,3)b�E��r�Zv�#��rH��܆fh,�7ή�@���f��=�f�K�Gj9�	Њ����C�en �+���)���;i-��q���~n��Y�e�����dF.a��H~��S�y� �]$�=4�`���*����^�9��T���tKO���b<���T������W�ޣ�cD�ɯ��	9RZ8���ZN�h�V��#Р��Mv��nL�L���J�8��sP?�,]K+
�I�M��wq�檄���e D�R����:��<p	W(�XQe�'u|b��o���L��gP�Ea�}ey��m�މD"o��hM���\\B�8�m�<%ߣoݫr��?B�* {��f������Éh�n:�Z�K�ș`ʬP*}~P�P�E��a�2s'��S�ʔ��/w''�/3�uː������.W5Ź���֞���w���/ʧ��%�Ɠ�r	�?q��V#��E�k��w�HU������#>�Hk�3Y?~{p�,Ld��w�*n2�`5W"	#^hLI��~/H��<�bZC^�+��Ԗ�	��	[/{Vy���[�,�\#˴�WdK^}�7��=k���U��*���bO��J?���6���l�a{6����6����'�§��Ƅv�d�Ϯܱ��޸q�	��co~�˵�v��S\�jc�Y|=?(��Q��m�S)a�A�v�)t߽���z9�b�"�	�ˍ����,�g��\���  4~�j��2ZI
H�"�{ �����uk��e��Yqy��1�h�F�3i�]�7걖W�Z۠�E@��s;; ��Z�����:��wG����b�}�<�̋BJ�K�N�
"GJ� 0Vf�yOb��J���hK�$.��=.4<�oYPjQ*~&�L� �A�6b��я_�&�e����L(����s��T� �A��ٱ<�[mp���@I��f�p�}kŘK��u�mWm�m2U����4�?v;�iE3`�Zp��e�J���H-T�7$ZPM����m�&�������X�6���3�����*7h�