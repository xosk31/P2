XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��I�� '��Z���T���3��!��h}
_��2A՝�q�F�W��;�R��b+����[�PvE�6}t��o��c�/f1}�{�)�B�� ��U>q>��(���C,���F�]t��'�����r�\X��m�Ў*��e~{�G���l���A3B��%�g�'�u�4������f�Wj�������Ir��v������������a�W@�������k�U4��U�����-���-]���Cz�dG�>�Ï���ef�-��eoB���=��!��;əj\�GM��S���d��R��S|u��:������>EҼ�+S�Hba9]��������hIwN�)�� �S��p^�N�4�
ƞkꢚ���sq� ����Fn��>�Q|�}�6TjX )���s�+<F�I}�9��!y\S�SLmڃ[�?r�Ί@@Jm����I L��@�Ǳb�S<z@�n�������2S�>���}��&�K��`&�:=�:N�I�1��j1��� ���
��^�K�°�Kڡj������;8�����ϔna��Ȩ���I4���l��Q�w�r���f�0� '`��Œg{ᨕ0(���)�5��o��<�!$I[����P��Xh_��t��X(_��~f�q)�)b��Y�$
�t~��Z�����GGU�Y����%�Xg��;�ӆF�z��ZQ�sD3�)�& 0B�7��P?1f��n�hP)�AxOH�@mTq�X��+����#Z��`ը����\}XlxVHYEB    38e2     fb0�	}���W�%��8���IVPΆ��Ǎ_�����j�<徉!??u����O�x����J�i���aed�Wе�6����AjӴ��#�͒f��TÝ�.��PM� �5G��u�ɞ��*�7�:Vz��b��Pݭ�7�'(p��3 ��Rw�k!�n��N�vh�Pqo�!l�bܣ����t9{�9'ɟ��%�h<����`���vc�Xf9�������<�OL���Ra��D̍cqR����O;��N���+�;�K�;7�U�䨗�;�I�������=k�����6*oS���9��8�3��߯1�������xkI�^�.�����l�fK��SOEf|��!e�wC%L��}�j$�)T��QJ��ۘ�/�ʌX�����Ј�0��eA2'	�AѦi��Y X�'nx�4�"��z	�SFUedqUF̶��/�r8{�#�z�;X7׮t{�罨�w�ā�p햡 �4�S�I�
��˝e�+d���jq�Q�'�b�s���	5��Ȗ�Ct�������b��&��x��wJR��-���Țɕ$ܵ�sQw�zwT�O"2��3�,E�R��K07�T���������ڡ��b����!��/����4E���"�VE5$s����-[�qp\�8�h��8�³����(��Q�bb���n�Е͍�'��"�>8�����V�Æ��y�����.Z��WD�`}�$9�'�<<�ⴭ�3&K�$�U�D�!�P��	 f]؉7���o8�ܲ"u�8y�k��{�����ΞS>=���[�վ�Q[KX���^{#�%n��:���T]�r������׃��.�,e_��,�Di40F�2_fOit=�����Q��}� ��ҏ�>���sG3T��O䟑n�3�ˆ�0�����1V��;=y�`�x^�B�7msq@z��X}�J�1��K�S�Ƽd�q�)?�9ԍ3k���ϼ6�2��C\>�_~��h��X3j���Iy�:�:�&���,e����_	Dޒ<#�ov�>>��]� Cu'�gCZ�}2*�.3j1Fٵ!�+Gp\O&�}�ѹ����$949-��-SdE�`�Mً�l��bD��U�g�b�f,��	0�w��6�E4�)�:-����pQa0�"��\��S��_dC�gV�����E(4kI�9���e��yC���~c����~�7�ŧ�{C
Z[\|.��]���޾6:oϑ�� j�P��y\�&���@��9 ���.�U�_zg���{��$�pz��N���&�[";��T���(�����o�׵-w��҈�{�[S��'� �I'�Z��52�F�SD����T��j3Q!�g)6�d�3�2�����ܩ`Ǫ;��� ���#P�?VfDP NN��#$t��bGؿ'=��s����Cs#��|�q���nU��~���3=Յ�{FR��:����{F�׵9@�-�P\�K,��C�h8}߲������ ��~7�<�e�[�ˢ	s&.9���	ej͟�Ԃy� |�~zhu^�8�9m�k�EB�����C��Q�R���n. Uo}rb;��5��Vc�}�Oe$a��Q�cU�{GVs�H5�����{qrR��H񂱾)R�
���5nKx
4%Oۅ>�5ʏ��iQy�Q�Y���H��fDT�����,���z��)�h��7�c©�P	l���O�~�����W����
���7���]����S��g�������x%�h��k<��ԕlC=��$�$CC��.���r)��~�ktf/��o�|4n(��7�NZ�&'-�T =�!^v�G{k#��^������E��g���pP彘�="
�����Y֜yeB���#)ԣ�b �_TvG�H�V0���<�ݻz$��Ҹ8?C��������+bV{"�����9�R���<� ��L��3�#Uwc�̈́j�����h �h����4Zj��$��P��6s�C@{��**�ɕ�fk��,�b���$����ΰy��l0V��;��,����YF�]��%�ۈ�Uiǯ�i���֭�'j˷��}���t
�.�E��|����>�#���6@��´.��}]�,�u�x̮���kS�"!J�F��?#9a,d/�P;?
vܶ�Z]p�W�e,�	�h���� <nM�%_I=��.�k�kyr)|��zѳi�^3̞Ƕ	��oY?��)Π���n�Ȝl����t��ʓ��(di��i�=��Y�Wfr����.�r����FF�+��4��ʱ�/b� ��D���-c�~zr��yo}����a=ua��	�H`�(�F�y6P���*Uk������[���K{�х���/�k���3#����Z���b6��>��I��eӈ�Qb4%��J����o��H���<{#)]{?�өpC��r��o���EdiFTݺ��n�M4ɏa��<�ڑ���+G?VZ��V���8Z6�����(�!��ՠ[gu,�1�h/Չ�f�Z��mS9d���Q�� e�m���6ם#�[}�����11bg�z҇�:`�r��*��y�lݤfmx��ɑ�ۭ����BS��ǁ��!e%�� �x(��M��GFUq�P�V����	(��X;SK�S.N�u�NZH'����'�)���gSz�l͞^��M�� �53�夯����ߋ�MJ0v��U�-��gs)��|�<�H� d��J��v��y�G��k �⾧�ף'ċ9�@� �&O�����M��SK�F:�Ϸ��=��Dy��pc�xg��; �ZP)q�O&�9ZZH��	�Th���R0�u�͋%0�*_�&}Q��	|U�����6����$�����X/I��U�T�y��_f0;�[8v����X���!�ZV�V�(�Gѕ�CB�>����rs�0�,?����H��XU�Z�6��L��m�+��Eˌ~�%�@h�3>ԪN�
vS�4��Ż�OMc�\'W͜�Wi�K����)�yaH���tpٓ�@U��0�R쒰�ꊠ�O�>��l��}��L�u�B
<�E�l������2�����V�<��w���2q1��i�7/��=��h�������k�Vm�*��d��ɧ�0`�ن��'@�i:xђ.�Г��c!6�Ʌó����!�S<�r�ź$L��tZ�F"��i[��L5��c�����a`��M\T�# ?���S,��1�E�{\����y ��j>1y9u���˦��_:(�R����*���k\�Mh>��a)k��Tm����������v�Lۣ�"�M���A»��rX�WF�$��0���7�,N(,�nW<�,G@��M�C<�;0�BM�� ���FC�Dj��֢u��!����h���f��a��O���X�i~변�4�$v-��4]o�aVz�(��e����H�18q��__́�w#�P���2���%H�3xۃA����aN�Q�w�{p�x�>�N�T�	h�jX��A�L��:;����W�����_L%����݆�>����\7� LT�qy���+m<��.G�:��|��0��ؠ���?u���;L�*xb$�9
=O����U�F�2y�R%;V�g V�0ьj�J3d�m;�+m�N�K@��M�n�*����R��u�d��D]�Ʈ�ө���:� �4��1�q���CNb��U�Dcs�֑o:��IE�m�A�V�hwx�ָK^����A{�#�;lcT��ox�V�:��ZZ��Y���NmR� �P�p}�&��d�҆$�0����-P��f������g��$�R�!yճ jI��D�����}�*pԟ�"��E�V`� �;�C��{]�F�y�"�eKGa�`��9��G�ǚ��^�eTGg�Q}��!�d(�ZA��8x�i �YǖG�@���