XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��1(�SМ'�v�,}��V���`�	��$Y����I����;�)��_�y�PU[q�/�L���r{S�M�f`64F6 x�m:�|$Ē,� ���⾝���@,��n�H:/X7�=obg�Jo0$���p�9}n��.P$*F�7�s�r��P�@6�1w��Kp˃��^I�K߿�Lf�s�1F��7-�6�w�k�E��q'K$�$pX������>T���Z��7BnOHɥ�ȱ֡��&cG��LV������e�7�E%Ie-�%��ax[��@]4?�ZrvC�{�8ط��p����#5��r uJ��Ť�Y�8(���cq:ѴN��s�ZM���PR�1����`��
��}�3pIL.cY�G�0��V���J,��zqC���?�B��}e:��ue�9��*c�1R6�����B�ew1R�l��{���P����7�Z�0�\Q͌�
�m123Z���w��<���� ;X��To�tȇm�����"��O�e-����!;����r�L�Tfp���Q�e�k{��|�!&��۹�+]���}�?�m:�L�F_�]d)�����L����+;�h(��4|�A ~!��8^ �:|5eD�S܍�����`�\�Ija��_Nc��$;�^.2>DV^kN<p�~ⶺ�\��>��0� ��9[�7I�R$/voi�D�D�1�_���!�_
Vg�j�kd �Bl�B״&���N���M  !C����I����8{�Զ�XlxVHYEB    248e     9f0(b�\��=��=�]m��yTc2[��ͫ����xkO�x��	в��������@H���/
�g�X�~�Rd�=P�qG�9�	Dӑ5f�7�c��%��~�$a* 0�ҩ��Q��҄h@"��w�#`�^�Tz�$�M��U��_#g��aRTƽ�F!�,ӉR%K��h
b����&�5�1��D`�<��
�ڤ|�U]�^��������+�R.��	0E:��2�[����R!Y�+���l��-�X��k�]|�G#��N���Sb��������;�Q@�ܫ��c�U�B� �Q�u^�;�����0)���'��rhB!i{�c���w��Q��`���V^kbG� S"v��'�m���0Oɿ�s����u���5{�{�wL�Z��VZ���Y�cU7$G��1R�4�L�ˏ������D�I�v+���0��!O4M)2�{��,g��a�$���q�Ʋ���Z���`�x�J���_\���_J�MS|��DT�4<'`�cJ{=m�[zBť������i�}a�z5�����\�08Ew��r:�o���6�2塲�-�֜5�e�j.G�h�N�Q��C\<�K��P>��IQ+��U׊���8�D���6�k9�o��������j�^�Y�p.�t��%��4ku0��Y�mb� �畸��9�����Óm�-iAݼU�۱i�(�S�R;�4��A�ɘ�s��<�	�W��ш9��|�\^4����S-��\��C�V���ߺ�*}_��Ť;rn�*6�]��y��gu,�zf����vw^�8R(�C0�4��B ��ҁ�B쌓�b��GB�{�����~9���w���&��H���ɵ��,�?�j`�Cl�&k�l�
 *"��3)�Ԇ�	���ڞ�I49�ׂ�M�C�_�s?m���^�[Dt;���5NA�6 Lۥ�,���KE�0�όmޞo��ZG=!���]^��a�E�w���֨&�py.p3�)��-$朢�=�
<����j�}�ڻ<cC����2�v�����6��!����l�,��A1�Hj9!k��9Yi�a�d.�����ox��! R9]�t��J��A�xD�ཌྷ&���o	8�Z�E�����I��ڗx��i<Z�-���
��=í����0����^��E� �o�e�Τ"���<��u&��j�-��8�ӈ����-�9����t��,{�xd�M� �Ypn��{��"��.y����A��؆��l���ŗ^���:Q�
��,v���p����N
�0|9���o�n}��Ao�Zo���e�AV�%�1�u=���/\-���Б��||f;�m�u̽ �V]�ִ���wD�S�T��#��pI[�Xq�����I�#ig����8v�W	�@�8<h�o3"�v����m��T[���y�y�-5�FԷL���F��Ќ�� �Չ�B-����e�q���|�Q�.؝dL�r(��i�_�B�Z����h���=�P��������� �}���[���� /^�ї�p��B?�I�(�t<Gg��7��P&�Mp{|6����������� ��}Uy�j�!�St�47g����8qKh�������%2���=�^�f� ��O�?~�+�r����㯄[�i����Gm߄<:����]�+��)Q��T�&�&���z+_��1�ʖ����ó�)���LJ!G�Y��?*��K��4�p�N׭/��'��oQ�������:��2`5~��8-��WC��!ɂ!o��k���Ϻ:�uc ��=���;�h���aC$W6 ��[��\�m�%��m^ �;��d���X�u��o����(u2MpGy<nt� O���\����&��ȼ�rڃ�v)w���vSi|����4����uPP[�vᵶd?����A1Eޠ�(^W(�_�ݚ%�u,gz��@�Z�Sf�dX}�<aWB�$��%����?Aݒz�m	�8�ڱ))���Ѭ�H��c��;S��H�)X�O`N=���*O��LJ���հ�a�Jx���sh�5]����!>�p.r[��Ş�E0�'���vst�6gd~@(�N��p^y���A��{՛��Ҫ/�������/4�o����(�T"*XH3������,0�P�G�B��j���Y�pO��|s0I�g��71���M郇�g���B�-ޟ
K�툔:`?;z�9Ҹ��	#���0��M+��k��"@$��u3���fL���b,��������o�VNjXǈ`L䓁���
����m��PƖ/�o��0lg^ی̍����.�l�j��'c�=XqߎP�_ࡣ,]��/Md��8t������:U���!��ѶG�P�n���n��hB���$�l,�=s���t&��~�𩜔��g���D���$��f��]�[Z-Ѹ�"�nM��ǋF$"MW<#A�VF�B=�g/�p�Q�r˙��n����r��Aȷ�kR��y.�r�N.�Q�&�I��c"n�ܾ|E>�