XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��W�O��ur�8�$����YN��IQ���)n�0~��@�֥���heķ?�J
1;w��_�/���w����+����a�G���o�u�}�Ԑ�?��Cc.�"����1@��0��Ř����(-?��V
n���Q�m��g��}�߳�����X{��~��ptuULK��Ico:d�)���5Y�n+��'�>/�(oYX��y1��Si��^{1	`��&������#�>���Jؤe�
�Z$�8�������ʨ.R�jZ��y{:�r�I���P�=��ר_����Z/��6a"�M���R�\~��LL���1Ʒ	'�fq�H�t�R],Y�:6;�/0VOoխWD��"ʣa6j��{��VM���������T��{qS22j3Y~��q���[�b��BB��':�J��G���ӗ6��j�J|��#-���kN;[�b�����/W'-�$�8�,�����px,��h)����j�8��T�4�H͵�b��}�`*6u�ɂ>��`ai� l���Y��C06��jT�0&�1��yi�h�u�x��U쨘�D�(�n���&ۍ��T]V���7RG �䏑��'���ݲD��iC����V�p�3ɦ�I)�Gx�2�[����]�l_�W1z�W�$7�I�t%���wVk'��$�.�v����v�]M������L���3;^�'�2��)y�T	�|������P؄�pʩk��c<������q�n��r�y$�J�	���ڸ�XlxVHYEB    67d5    1150kC��(�t%ه��`;�?Y�,N�A��Y�J�ʦ~J6�6����L~��/\)FZW�4���\t���r^G1X��/�U�=�����J1�]O�
HGL��߅}�.�����c�#���.ZV�p���ϱk9)�Ұ��-PC8���؟�����xጨ
:*�uY4�u��1S ��o�� �(�4�.EM����@��*k��X��~}B���i��-���Ղ\�D�.څ2{���_V�iN	E4�K�X�|�pͦ��yޓ��b3�S���Ѻ�6X+�̸�з�q�VeQe嬈1�݄��iޓe���I�s��r�#����t��z�Tݷ^x���_阑H��W0��kP������-���׷b��X&`�Lv_v�E��{�^?�/�a�����L�����z$8޼�
d䟊��}& �B�#-ᨀ����4/*�"�DT�}��/���
fX��x|ζG�pCb����q&S`����Z@eJ/��Řu.��,>�X*������T;��?Σ�h�䔻K��y����Hxbi�)B>3��)�gAt� ,�򺲜�l0,Nǹ�h��k�E���C߫Eq� ��B��}��]6{��v�TB&K[?j�<Q�V���f�Ҧ(��H�r+��O�f8�x�������-s���s�`L�� �:�WQA�qR�k!�55��} b{�c@�m��������Ӎc��T�O5�ͳ�c�/|�n'9<��㣛µ@,o3<i-���C�3�����͞����X���~/�J;7�?�$�ਛ3�����7�6������ԋ�6'��n7D]X����G�:{;��Mj���?��vPG'�mf�+��O�ɉݸ�L�.�W)q�\b3���7����̀J��������������nj@R��v��Ǯ��*b�g<����\����W��jR��L;g7��T�U$C������8`�2�p��.�P[���j�&�T��(#�L�M�s�"i�!������wA ���k%v�yl򩹍+�=�Y-���w�.<��Vr�%�5�up�b�h0��]��֩:,�g]޼�Ԟww��t"��
�<�nW�!�ʹV�����٩�x"��,f�(��0׺(%�8,��rgw"(ZNw*B
��\<���l��	jK���7ߩ�Ēb�dwa�w���)�ͼ�Y"��)W�rq�'ύ�8���i#�B��D��S�;�O׎�$�)��Q6��$-(��\0�m�� X�<��c�ٵ�<�����!����|#��2[���-�r�ᮿ]�7��G��7��	���f���3dO6JB;]I���j��<�u�WG~�����#�[4�d�N�s	~���빰m^A�*!���O�M�$n������Yi'�O��~�R'��8#/k־7J�^G�q���w�ȎI8�#&�[{�j��'�ZԴ>�����:�T�L�޴,dG�}���[F�%es��OhV�ӷ[m�r#/Q���l3�L�����~%���"7 K�;�<;�XCr/�/L2��+��e�� ]����꼦�s��6�#�+�
�����^��02����6��/Ъq���q��:.�~_�
S��%�Mok��ͨV�:"IvCy��k�-܍��� ��M�K2v��U�Fv�y���ᤳ�:!�?>, �Nw����]�|��Dщ���Ыob��8�,#)hlQڭ�h�Ӥo�g�7�������+Jw��f��'W��}Z9�>���mA@~-b���C���kІ1�Jѥ�L�T����|�@j"�,�P<�-���+W@�f.�m�L�b��9�Q�{�[��%&�B]�2g0;q���d�'��MXs�[��wp4��f��zd^�}��I;��t˝q$�����(�a (iԂ'\��J�0�b$�U�& ��%����	?M
+����8]�$��p�%V�#�E�U]�C���l^����pH���	ԁ�aIy��d�iüY��h.M���R<k���xYX�ǯx~l���`�w���Ϗx�_A���5kj��O�+FH�@�^�4/AC,��r΍�b���X���I��v��Y
����am���`!K]���pۂ[�̀�7��b����w�0�N��5g�Ӆ�]�gKA�pU�L����!~���f��~����8��-r�5����@"���̹�G����XW���wSQnoʋY%�I�s7755����W��,NB��YO	 � >>6���Re*iZ��f�w4��*��P���~����\���v�+�$[��{Ӕ�-�W�ؠ���z���� �3@�]^G:���g*�S�q��^��� ��4m1��]�R�C����tx�Vh�����"(}���G ��<%��c���f�������0X#�x���%����#e
O�A��<G"r��ꩪ ��o�ʶ��
p#g���z���Ā�Up#���/뿦"Z,�1�T�k^�6R<qz�s�s{ns��,�U��0$��3� �l� Vn����*������(�X;c���� I"�%v	�D8�p�C�Z���؅�hrU��������??�/�%)�ј�t[�R�%��F�C|ճ���f8H��[��"��	���ۘ�V �����;�y��y���1(���o,�y7R������3+���k��l�^r�*Ll)+�/����C��`y�7��N�ŵ�D:��������[|�X�����	ģ���Td7[`��1�q�#��*�q�m����k�Ne�?�(֘�"&�]��n��8�>Mz}�YG�4�S�~͂J�d�,�g�� eCb8�t�_��[����E)�>�=�?��*�Ơt���z7
w��s-�kG�S<�����!�ȶ�t�\�>CP�I����rw3�0eǌ;�n�C����4oV�zX\F�Y�j^Js�\��9N(��Z�:�1Q��WZe�����e��,Cͅ��L�Dh/�Ysg�^�Rf��k�*�nE0Fl4��H_�{I.��Za��S����j�2�����q���c��j�y޺Ӄe�~�@�su4����/E�]~
��FUq��{�8��9�Z�l3�ta�ف��%S�ǿmUaϑY�?H)�������"�f��̄GS���+�
8S��f�������?��/����
j��v6?�M�;*��@��;w^E�zȹ:����X���R֚):H�����Hy�����6sqػs��?���X�="��t�t�Y�[ݍ B�&[!�ٱ_?X�� ����y��;�4����i��̹g�E��!s{e>��]Iu���D�`�gCY���|��5��!�c}�S1Ɉ�Xx
�i�._C2�ľ��0o����j���]V���0�kf�q��T{����^>fP�	k�R<���*w����!�s�$Oa�nKi�8���'2�ZM7�v�^j�:҃]������vT���QeOV�;�����c�Gp�������-�[%�cZ��r�9�c�������'�V���Bn�:���s��?�_?���\wu����%�K�#1��1�L�x~	�,���Dq�{:ϫ]u�-&�?�f���s�Ŝ]��Gk�q�!��*��7�@��^������0����-lܾ7ؘ]��3����trp��9����?o�6Yn�?>(�zZbt	����xN�̴��,R�-�1Y��&��Ʉ�ڸc����p�?���x����pqӌ\
�tR,���f�g��4 ����ˌ̦%�g>b�G� /[o !Q�i�@9����u�D�(�9y��ϧ���1��MTd��:�[��a)w������3���!�h�5����V�D���r��>��Z��!�'"�/I�]�'h�Cߍ��y��F���0u�8K���_��R7!�
I�%�o��̱��d�3\W���U���3��Xk��\[�l�b�E��|v��۬���<q}�R��;��q9�����C�7��k���s,Ou�Ɨ�
��=����ݚV@���7
��0�f��ˁ��[6��i�V=�ڟ��;��Q	i�ƍ�뢢fA� 2�<���uKM�F��W9��S�b7��.�V�C1��RC�@y1��R�A�S8����@>{�%�%������@ZOl&3��fK�_����z�� �↉�"��&�F���("��ʯ�;V�E5���/��vA�6�{o�2�PA��?p����n�*TN�C�2-��ߕ�s�#ϐ�8Oq�� ՊT��X/�m�r��Ҥ
�.J�=L�d���.T��XH6��p��ԏeZ�4T�)i��pL�@