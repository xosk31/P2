XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���u��%���X�4u���X��[Z�����������0==�����|�t�rBJ7�Z�x��P�$�r�vƞ�a
^wt�� )pǛ�M1� ���T��ƣm|�ʶ�J�k�~�������ϡ��j�x"9)C_�r��]|�<V����ȎHLm>�����z��5%�H)���;��I�3_!��:~!�(UH4���:�!ia8@<��r�1ܻy�G���5��ƃ�ve2�@d�H�x�n|���eۺ�N5:�
(���
=�a]��qD��0���r�c�Dm(�Ҥ�xӮ1;�ߗ^��6[A~�W�}ʬ��;�����P ��x���ek���i����f��
����m]E	�GR��ɷ��X���]�qA:�'�թ�1E&i1���v~��C�Ϻl��r��ӵ��,�4�i��)T�m�E�%��Ĥ�M'�!h^>&1#���"��)�+t LV����)�R�?ǔ�81iW9	̲��A+y��B�#�6���;��m�lc0iNƮ�gB(̤|���+�ia��u�/��}��������V�ݱ���*��a��7��_�����\߱hh���-��������]m|�Ik��r���,��$�#�Ċf��|ؓ�%}S��7Z/�v���Я$ʈ��}��"���Ϧ{O^@;UO�� �����LW�\��ک�壦�� L�R���S�뇋���$x�P�e��~�T0��5� �%�zA����6p#�qXlxVHYEB    c3e8    1d20���|�����X>2e\=ą��Eۚ�Y��ʝ5�ƭ���)�:x�}"$��~"���
��Z�{�o�I��i�&fji. ������}�z��V�(�ћr�ȼ�;zgB1�G�p�*6�Z�����Ӟi,�},)XY��/�@�:b	��^�	�x��$֍��e��#��5�6�5�T0��C8ػ&�h��\��3��|$�O��<��y����(=�S笏O�*z�z��V%���J��Y�GנA���co��5f��~ҝ��}�T�~�����ߩ�U��>�i�~��
f���	8#��\sG�A��.�������5�����b���ӢVeY�^���4?��
{F�kk���W����pz$.�sKu���?��)#�#f`y(G��lz�k$|K,��IR2d���G���]���H����<���~¦�b-˱����_�K�B.*mz�$�"fz�4���S��OT�[�B��Q�]�.$��IKvV��+}�sRU���B�"�	�׋4.�GRPFfCܝ]]��#�X����gퟘ�z�ے"�7]�
a�1اC��'E$+ͳ��[�Hj>-st.q��Pͬ��P�%��&���QNW��p:^�q�:���G�igfy=))h�~��l10�Z�%�[n� ú�����ܐ���v0��1B�2��0�b�z;*��6��'$/Fܩ�ae�:�crX:mY�� ������r��l��qh4�pſ�$�Js��ĪJ��č�өgVT��Q3��s��W��=f ;:�������k��]�C�~@���Dc��B4��T@�!8(Ԋ������R�]$Zlԭ��~lF�� b��L2lW4��P����H�+Uy2������w��0��~��+�	�������D����9�p�Rs$k�4oۇ�ͫ���wA��?�Q�E��2��8Β&�i������yb���EI4�a�ʢ@�eW�Ϸ��l_�P*GX��Y���V	�P>���;��̓K6B�XD/9�C	����M쇹r�|?�4���r؉[/f����i�����,��V���
����gj��g���j�c�|-�\��[�3yH�XQ	`�\5+.��U��v�J���)��/��a����)�7��b3��V�^�\;TO)y����Q\h�}��C>�RO_�A7�	�6
�L_�ޟ�3�+�I��� *E��V|jB(ȍB+�2�j�r�eItM���+��R����<�X}����Jf7���J"Bɝ����ߏ�h�L�0���#���~��'�z���jU�:K��ɕ�_�Ip���d��,��TugOM��鴪���j����D���m[ZAe�C���=#�O�0'�6I�"Y[9�L��9~0��}�">(��Zʄ��ە�T��f(L��{1�)W�O\�_Z�V���"�!����Ƴ#+]nr���[}A�(��G�NN~i	��Y�-m���J�[他�_�'��BtWQ>�O:᳛Rv9����v4r�s��r�^v. H�$�`vv[�<��F�ԑn��YH�����x���cʍ�Qo���ƺ�����G$F}D�Ȫuk�<%�9����U�%��,a����b���r~��r���������H��ҧ�`�pJ����v�$�q�?{Cb�8�Oss�<Ba��bb:�E|������H�YҢIh������l�c+,������X�@�I|��*���ʝ�]����I�q�(�!L���j�cc7:vQf��<�C��e�J�4U���b7ř��d�%%���E�F���Y�Ձ�m�;D|�&~�����2�&��5L\�9�J��H�X:��(=�$m��*d���>n�;����O����R ����l�Y@��9�b{#��C3T�Ja>n�����1��I�6��s\"�|�!��nq�(�`�7؛�w�;���	���o2�+�u�"{F�q	;.o���b^kL�������7�a/��b�!����C�9�R� D[����;�5����i��Z]�&H{Z(F?Cn��j��?�f��wI�:~E)$�J��`d�VTذr &�Yv8�bF`����~���5�	��*rj�<�6��CE�i�E�O�IH���(�<N��$l*;|��k�^�}����m�vNUD����Vx��i�٢�b��&FڕHMęk�
�]fz��'���/,��59C�� [d�u'��}�� J78��D,�'y�Ӧ����Q;�ƨ�����&���,"G�S�q!���Bi��4k��b�����XH<�F�ȥ.}��Z�O�mP�	�ꨓ�Ƥ�X
T�ﺆ����J�c_A�����d��alay0VB��6�7��E�e�i��kek1�W�O.l�Qz�
^�o&�?O�F��(�՘+��d��b�zU���I�CL��p�����GJ�t�]�8�E��d4��Im���`빸��2WM�)������}��_$yP���(7-J�²? _�3c3ӫQ��A��6K�X������2�!-�-2m4�	�dʵ�������Mݝ�[���_�Ҹ-��ѭOW��o��q���#�A�>S-�"�`u;����ȅ�f��Y�`��9Iw@>5R�C��MzKqЍ�@��olC��sη�, H]�C�h���bb��a�y�O�[F��{T��@�[t���ztƣ���U���59J��XZ)O�e,����w�vK�%=�yJ����!��7J��il���u��� '��Is�^�������gQ�H�HU3�'���><������+m%�V�9�8v���3d�ϥ��n�ގ2+�Ѕ����t_U'P��C��r�ΉK�)��7���ml�q�bh����wt�p�L��f4
��G�� ;��9�u�oTC�(ȶg'=}.~<���?[����̮�Cǿ����p�Ld��-��S]=]}A�8�<#��]�nn�}Ж�Ó�PZ�*����'��؎�����>x�JT��{�����z�	���Fz�'����`���O����w����[0�	Dp5WNT$�����&<�:nk��tQ$���bH�p�иռ�����
�o˲g�8U��d����v>��/)�LU�������}u��.��D�YͯF9OSs���x�y�j�ug�썱��X�a_�(��Ώ��{��K;$ކd�8�4;a�� ��ʶq�8�λ���M�6�$鿨�׬��]3�����i� ���x$�F��R>��8����3c��f����1�Q>��w�!�nS0��j2�-ބh����H�qp���a���H��=
z���¤�[�RTT��7f�	�~F4&?�A[e��`��^�tE�Ml���Y|�Z1��F�B�	=l8�z�m��_�葎Ze�|O�;&LLJR	y%����Z4#���n&�AS��P��.�#�W�Sh�TS�w�m�=�e��dW;�z�$�Y��s�
��h�=)ε��A��t(�d�A6���d�s������$x&΀#d���$�&B(g5}~b*�nN���OĬ�/v����k��b�.��O��_���y�*�Sa��?�S���l�%댳F?��m.�OO`�y "��0s��&M�D_9
^@��k��̽��ր|�G��r#���E�4e�]L��0q�u"��<�w��۞��b��si�0�k]�S��̙���c;^}S�T���q^!1�T<@ߜ�(�V7�p�$iR>��u4�k�?M�}s�:�*R/v<�L~����8���ݽ&i�������/`��C��[��f#��^����Z�7��W$nOdi2��G���f�٤�8/]a��.�r?pZ@}�}��4��f�bd.��;�uK�ƐDcmu��������_�rz�o�'��`\����w��BZ��.)_V�Lז�a͏Щ����r��������f�m)��kO���L�͙~_�gS�jB�Ģ>5���;�S��'Lق��ޞ�w��bݿL(ò+Ṛ��_=����^/R�{	���+^�B��_lzR�f�$U��w"}ET�$���>V;���y2�����1�^
���ǔ�:v��B�J�7v]j�2y*����~�rV�4B \��W� �+����� ��2���s����� ��8��d*w�O���戻���p�ڙx��Z5��;ڌ���b������B�e����e��y`�<�"F�쮢~��i@���)�v���bJV�Y�_����?�ȇ�)v��\�^S�g�C��ہҎ��>1���(�8t�Κ{a��3���|�s��j@x�����z�Ƞq���D動a�;���V�b|"4�FA�c�Ai$#�pJ�چ*/(�����v=Tun4K�[$d3a�'|!S����S,O1t�=@w�s�}%H$�x+8��Tӕ�X�����M8{ Ț{�d�	XQ��a��4��IIE���wg��H�n�əo}$#,�di�Ѣ*����Z��H�0o�Ygy^��#b�O�^8��{�6�G��9��<�Qa���C��õ�ld��v||�`����sŬ_�Mb��SQZLɮѣ��Z�;טT��i�����M�"��`�e%���QP���6!C�$�J-�wS4�J� ����9Y��-�����p#G���_O�=���*�R���_/��	����w���^>���ؔ�A'�����YZY���c<�pg��5ry� ���2('�����0��5�[L�D�S7��s���I�Q;�����P�SɅ͑�TBF�ԡG�����H�4��(O�]��85��>��n�Z����w_ ���"xR���[��g��r�����6!	埞��\��x��C�bk��V�1j6��De���0d�+q�Fi_�y�W�˷�\3�S	��B����[O��n���5e��+�v�̻�!hI�I�%���"�q�V�nf��^!�<݇J�
+�z�0w6a�E�ٯ6>�&ʯ4��\d4>�θ�1�|�����\��I:���Ud���T��a��qޘ���>�gW#��KwB��ʲkɕ1&{��IM|�5�J*�1�����5�/ �У��i�u^��T�p&+N��W�3����F5݋�@���`�a�.��Eʪ�pc_�d6��/�e�/xx�Ʃ[?�������>	��I�[�Fd�O�Z&�{h�񛧇ߖ��~'?O�+��/�r�Qb�E-F��X��{~D�6LT[1I7�\Z��}�R�s�v%�Z��e����@��%^O�n�*_$\���0Mמ[x�"�`�=J޵���0Uh2^���
hv �3�yVH��p ]�38a����V�7*�`gi����=������F���5�q�����kzHލ-��õ�t<t�/ލr{���k�\\����G��V�EߋgCZ@͟����f�H)�<	�")Ѵ��qK�߅�A��ԧ�a1� O�TN�G[#n�>�\�-|�r�j<�(��wj��~ˉǽ��B�F��#�TwY ����,2E�x�5_�T��$������b����Lb����y��f�"J^*eM���. V�Ȥ��D�����ǐf�1��=�O.ǧ�
�7U�.9�:�.}uP͍z%Q�Z��ז�o��w�*r��7�j�	�1`7�����K�Èe����c�8`6"�&�-S��]�!�e%��d+�_1����)�5;�n+����T
��<du����F�w
x����o����P�c����e���AI���w��Yd�k2�Fp.11��1��h1�T�'��SK�lRs��! ꕣ,(.�)~�W���1)Uk��<��W�w���y�UN].�T���JcR,,pB�u��Ч��o�yR�Ա �rz��BS�/F�ȋkS�	Z}`���h%{�E����F�t��x�ۑ<��L��D�h^W��L@R���.�	���[a��u�!�c�(�WγP�u�~�R�2�o��zH����.��	��G/��I2�
�%�ʱ|�U����f�ع�����߿G��t�WnOr�=��ב2�����'�sn�<*w��7���0��&ϟ+K�U�9��	�dX�Vј��Ө�0���.[W�]��0sMC����F�^�ݰ6o��-5,B-ozB�-9��J2k���_��}�@C��?��n�
��_�Ȯ1#a���t�#��^�Sj�-��'3�{��NvR�)�(�������o�>`8���X;� �qlR�٬�����.C��2R3ue�3WI�Jb,�7@���-�;<3��}��ej;��|A���Н?ʆ�Z��Z��]�G�תW��bh�ǉ���,.H����u|#���$C��-[7��z�[J�.v�!7@>�SI���Xf]�m�Y����2����3N�R��4�fW6����Q��Y?Vj����nߎDދ��a�C/H`fR��87v`���/�<��Df�|�{�Dm��յ[����d}/-Ƌ1��(,nh���f�8�%Ժ�`Q���x��e��+�Jj�C���������[.���iϷ�ov�e���珩BźLx���b��ޭV��R}��c�����"��+XXJ�h\kT���?�F�#���/l��}I=O�0����/�Y8�oL�Pj�D�x���2ʧ	��K��4�ɵנ�Ҷ���+����������&�ȯ��L��X&����L�ӌ�W�xH<�����Bb}~�t�a�?TW_�|ͅLE�6A.a���D��uC��A��?��I#��Z{�3yVhY3T&T�֌*��n+�N�U����b�`�c�b,rw6��-�V���:��"?�v�P�72��և��Xo6�O^h���t۞�|�5�!M^8��������u��;^v��֡����F�Ɲ�ds�qg��{�L��j�&r2�Qv�.v]��/�����eL�-�0"/@"�	�k��M9F4cKGEI��`3gֽ*MU�w�v�}gy�t�D=sB�����*Si��S���r��G@x�y�l�%�!��%�Vߛ���%�B�,�'��~�h�Q��BXCe�������*�����T����ۋ3��k�w����B��!�a%�4f�i{�ĊF4A�p�����#?�ZU49[�Ɲ�[d��Sr>������ǧF�5�R��ӆz�)���W���5܌��s(�{�"{,��7!G��RBNJ�d�`|T���q��;Ѳ�6*�iX��6D������M�,�,%F	��UNk2͠�ģ>�B��#���F���Q5�R+�˓�{aN����Q�