XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���d*n�=^mJ�j�e���+���<�r�]4�L�@yo4{4ԛ��FN���Q�+����%֔��Ƽ�!����bJ�{#v�n֥`r�q`��X�1�̆��?��l�|qq���h��`s����s��4?h�}�����M�gk�qh���Q���o6�QK�c(��75�����bd/
�!>����Ԩ�'���[s��v�F���E,;ؐ���^���G2:Z����h�d'Ɓ��X���g^It����r��p���9\�+����U zp;$���Q� �G̯���iK��õ���1{��[j��G	!�ɕy���k+��N�8:k�B�2H-��2Y^T4TI���m�i75{�<u���ʹt��@,Aj��~P����L �h��i�L_��M�v�6ӣh+p�gbX�[��w3������ݩ��*��t� }���ѱ�o;ʦ8�C����*�� Y�b��_�(��e텛��5�DJ�kW���N���Y�}��߫[L��O�`�r?�zz��G�	�\ r�е��k�&� ߗ͛�`'���^˫��Zz|�wz�L��pn��K(��bʪ�#+J2�Hv؏��֍�)dʯ�R����}��d�04�ʋO�hb�����政�o��=3�L�zG���ɐ|E����)�����퍏�%%�}���xy�B��%��?uW�ڳv��|-�\"��$��΢��\�"�Xqz�e�}ؠq6X�=Z�+��i��`;���� �[7XlxVHYEB    5e46    15303j������@�K#_r����/�{� �[lm��KcH3�P�e���	\ԃ	��q�U�����lۊR.ޒ,�G@�˪�&&�b{I0�G�g���f"y����m`�e�xw1�ɐ��.�_�>Y ǔ`���:�(��+#'?%ގx���h�$jR-(��y�X��G�	�*z�ߘy`�w0��+93�� ������4��R�;HE|���h(���1rA��z/`�f�Yeͳa�4��ؽ�	Tm�ÀN4����V,����d������`�qmtQ=@��;�Ǯ�0P�KvL�'�����Ѐ_���'�#v�V*xǝ.� ��.�T#�њ��<�g�(�n40W�8���l��]�b)\nO��w�7�e��|�4<jA��,�� ?�Cs�|@ԏ�)t�0O�ٰ�â_��څV�W�&uf�ʹvV�8AA�!}X.��v1�.�@��Ӡ����ě����yTr�YvŬ�p�F\���9,��	��GG�v�kpQ��e�o�QŅu�(q/�Z��
Peg~/�A�"G�ݻ���;`7�X�k���%'�/��VϗmG�M\H@b�ɉ�U'�ŽT8�KV{ �գf$�:��I�N��M���qX���Y�ڵ��D������s^J,v7��:�`�B�U�W�E&M
��ƥ�m�R���������.p��U��x7幃���s�Z<u&�{.+촁��]��.��je�y�X�iM�Xvl��u��`}�m� M���ڜ��? �꟞�zu�@�tn���d�"4����&�/�1���0����L)� �2�!!��Pr^~t�Wg�Y����(sQ+�v<�ܷ�I~��Q�xᰚ,n�q��eC�wP��9*��)��H�b`��K�W����'�`>a��f��.�AR ��T1Gw���N1/��N�
�.;��ߖu��EI.�Mq�?e-�
�M�۝�m��;NjY��(�JCSS�}^eێ�O��Fۼ�I8㰈0�Bλ�!rU�з���ҽ�T�.���'�U"3���r9�r��.����W�_��,.�H���Kt��!�����mkqJ`fu5j��l�i��Qj���)�:���̑��|�#��01�(��VQg�"�1�ݏ�Oy�g�~L	�vcۥ��N�i��;P�����q�A&��
��k��aŜ�2=!u!J�@4J�K�]jt��d�q5Q	?��ae+.QE�Tɟ�O�d�+\��ʛ���81�����"|�q��K�����̀ظi
us�k���L�+G���w��fiG���-Q�7�71������8���<B��)h!���K��`�0�ZE��HՋ���ި�)$/V��ǗC����N��~� ��D��Y��(H����kD�*i�.��b�RU���8��'4��p?i��W��r��h�ꆾ�;��x����	.۹��a�����7�����N8�Q^�Z��#�_��|���D�&�����h5s�ڱ��j�{�9ʍ�Z����`�f#o��|��Zxq���؈������[?Aa�|��k�5�ܧŶ� ��j@wX�a�+�T �Ō���^Y����^��sO��K��>E��ik�l��;�@�����<g?<�Y�N!��<�J��v2��L����))�:�c�*FX���6yڌ���Y�{?6rۙ����+vx,��3��0���I��/(=hݰ,�s
2Vn��^��r�D4�ýko-���y}F�k��{����,:�<=�*Ճ���}7�W�5;&U�$���l�!v��6(�?0���TS����X%���/1>�E��8�ޮ�-!�]ڧS���;�/�.��޵L��ݨ�x+w	��2}���N�<�U��8���}�mL�?�vo/���B ��������h~�+�p˄*��_w}X16_���zT���,|�}.5x�I����NA�@��v�mn�}�e.�]����l��C ���ȇ̡���o_�c�>�A��}W�����tk�����ګ<mc�-�;[�T��n��H��m�����x�	��j�+��OE�c���y�(x��TS�T(1�o	+Ś'ϙ74_�B{�&g:u�$�E��^ "��%k�A��y'٢Y|���?/>1�wQ`+�n�]4DnN�/����j-�� 2��s-\"�&g�,9ǚ͈�E��n)�`����_O�<�V:�{w�����Lʀ[�8̕�ĐS��=��>}t!�f���3+�7����L����� F���"�B<xfR��%N�ũ��K4lZiN(	c
JB;���������qR�Z0��YIך�ؔyH�}R��� R��w�̶�5���x�P��3CD�ʺ0��&E[���R�`O���[(��5�|������.N/G�T�J4�Y�f�PR5�N���q�G�\32�MW2��������f��)�;�tt�7]�TV�,ys:e���\-ʭ]��%1[��|��ԟ�&n�W��ɧ	L~��t�=��o&��S�6��(��U������#:��	n+#w���0xϲ�A-�=�e���N݊ٽ�6���V��g�U�{4���Y\aL�R�S������+���X��z��@ҫ�S6ic������~���W�oKqb���Z+�a����i9���^�4.W,���kzx�b��{���씽�x_�ǋ6:DmQúx�n�|mG�Ó��pl��0iEp�p�)$�� ô!g>��p��<�����Xl��k2���D�\��`�����q
�e�'2ˍ6�VDP4V1�]����v�F�N����-�Q�p��y��@�Q��U1 ��Za_5��guxP��7�E`�����[�@\��4��΢໰�D���ո�@f���L�u նN��h_)#M��b��)KJ�^x?ϝ"�C��c�$�hO�q�t�*X��+sfa;���r!�<��	�T1��݂4�n[�MU������oj��=�-]9r��_���9a�&��F��� ��`��*��U!`�_yxƷ�E���;�G�t�
��gF�x�⣚�A옖��������'���>I��[�%��˻�3�;5�/��6��{Ǖj����4�&�Z1�Z���v���;�d�N�շ��r�.͑�	0�8�҄��q��J�����>^q����3i��.����K,��]�L����7M�}q���vđ�(Y��xď��I����e={��N��0�-G*%k�޶Z�GL׈��WO���M	�s )*:OX�apU�L*�Z�~��Q��swcw�&�a�OȒ��	�@�g$��$@����]�?����J!�T.�)t�&u��D�bvcZ���~.l�-��d�A��(�1g�I�A#�+��9��L����8%�:@p|TDD��X�9����!�XjĠRUG����J���^{��j�ۯ��v?����{�I�����#Ӈ����<vx�,��cbs�ǔ""�o���`�.
�t��3Rv�Əa�/0��#i�v���N�q~�}������4���j$E�Z�W�i�תs���bC��sG%���{�L���!��h�C��i��{��QЛ��{3v�@pm��]���1<����*�K���7� �?+���o���6p	*$�ji♼��;R ��?R \"�t���vX�6���,�D�b�/͔��������d2��c����ҧr�$�K:YE'�Kzΰױ����h��a�'�����H��6�|~v$�T��-�o�^�.�yO�� $k����N�3A��x�iH�Ϻ�W� xJ}�!.B>:�@��dt!#y���=�^�@r�P����(C�E�+��E��;�t��$d�>>ڈv��D��,.�r��qd+7�	%�!(\��g�%�G�g����#|�8v��|�p�!1NG��DG>~p��a�`mt���{)�>\�:�>^ZVx�b�I��A�p� �������=��6�ȭ�9U_bK�Yƕe�Z,(�,�ן��<]�%� �[5����d���X�	A�?�La(wl̤��-xIh��?u:�_*WUd�f#C����bk�K�99�Ϻ�>2�&o�=w�5}�	ԣ� 
\�pky��-����P6���e��y_	U��3o���m Y��-=u�´�Cܟ@��퍁Ph���w��H�#���Q-n����F�ǘ�>ւI��V�=A�����f���
��!M0^�H�$�;�F�mLP�~�'������H�Z�c��)�����!� �Q� h|v��g�%�Gǜ�y`򠊱�k"�κ~����E�j�~}3;����o1Wl���GIZ�	QB�~c�f�
v6�lA�1mj�=�vj�q<K��T;��5f��� 0�M�����c$�_N-LO��\!�꣎Ɩ<�8�bY2w�g���Y'���Gfd�>њrɓ�������9�7.���E޳�3Ş}S�pq���-!���O�o͕y��:�J����6s��|5��W\��&71w"z�j ���2x!��.��>������M%<��5ŦK2��Wˢ�vcs�� Dx���z��ݴp�e���j9q�e�II~��x�Z�Ϗ.B�4S
ej��Ŧa��	����f���s����4;�� �	k�x�!w8n&.#������X�]���Ѣ&M�H:��BHHe6X��9�n��[iR
���j-��2�p�劬�F]���;����x�\v&z�b��V��?W�̭9���S6U�j�gcY�4�����;h׍�DшCwNx1�j}�$U`�,#���&�>�(+�E���3�a+��հ��T%�z9���3����7�$:kC�=)��x��o�Pbl�[���Z��XZ��a�&3y=�y�5����h��-{ ν�E��Qz��H�iW�	�D��_Q��D��Ro�ǻq\,M����7i}G���웋/~Jg☷�ŕ�vo����؊0�@�����ʊ�9�� 2
�Ɩd� ��O'6u7O�8/Q��"��ĝui��:>؇� ��l���M���FkF1�e����`��I�m���q���ɼ�Ýj���3��D����'��__���/®�~ �qy�*xI���(���2w��a�=&�i%!e* �̭ϒvV�Y���V��TAU�� Vf�=�_���\��d����a�`6Ղ�7��x��Og�]VD�pL5v��rD��Y���6{��n�'ͧHn�7w�J���=�x�˚�,:
4�ӯ����YΎ<m�9�/96���|Ɂq^d���e6�H@�����ű���G�����!b��jrCY��k�����ʉ�4X-�ܮO= Vb/��p\)ܫ��