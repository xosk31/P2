XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������t���Y�S���x�/�vs褙���Z1!�Y}@ĵ*��%��k�!q=�� d�e��_T?���a���^���uP&���#�=�#�7�&z�J�4�g4�i'�ue}���ˑ�S-9��g�\QS+�Nn�.���C�T�G��4���x����6n�?)�i���Ѣ�C�@��q�Z�j7�([y���X�E/�&��3�!^�n��?��E�]x�2�-:d��<D;��_�%j`�g��p��?[>�.��>!��$;xÔ��3_��,���ՠG}��7a����{W��Y��a�����#����-�M�\����.{��c�E�Q"��:mRD�|*�s	��v^��ͱ��_NP�՘��Q<��48�I?,��5�T��O[����94��^F�L��8'<p4�r�KR�������o�ܤSK�"��W2Էˤ��L�5�Ӏ���������&^q�S�$��d�^�>� B�}�i��AOTA3C�\Q��$vuv���'1�������J��<v(�}eJ����v>8�r�]�?�!7*g&��O�ڭ �2���#��f>���pV���#K�p��H.�ո!�>b)֖9XU0���P��p 	��w5g�n�q�����:���;�w�l�����1>� )L#sm�!B5�;ҩ�Ⱥ��t�]��*EU��+�����}T٢"�@K�ƹ)L���}/�	�XvC�2)�J)�b���R�>�#�&|��
���%�VG, 7�4��F?XlxVHYEB    4f43     f90,k���S�Һ��0�nO�ׅ���g/B�՝k@����z�VON���)� _�~����}�9�E�c���D���z�[-�Pnq�g�:H+��*���v�ռx��GgX�3�|=+�踲,�I�ş���ׁ�"ؖ�_�C00��G5iz����ꓳ��rw���8���s�����w�Zs�5|%<��:�{�>��k�G1q�]���}S����[65ʦ�4b��b<�W`4��B�����=6�|�����]3�n�֙�M�H��87!��@�q�1�,�E݃&;�wUk"�kƆ���B���A�E��57w��a���9kqެL[V�wg�^{��}u���c%�j�O1�G���]�Ef���|K#)2����Z�vY�����^N�6��dQԻD�L���c��R���v�9�RT�� �?�?Ee���]��k1P0u��'�����}���u�ũpd%zL#�v���c��f�n��e���<�'P�6&��Av�����eЊx pB���L�WѶe��,29�	/}�1+�s�9�ĸ�o?%ߟ���Õ!u+����i�!Ȉ�A�^��ظߜ&���{מ�˄��	���rY���O�3��T(�U�F���+�>��l6�+���a�G���O�����/�t�۱�3���iɷ����7�_��C�d��U:q���P� [�F����T�����C��!��|�D��M!�����U�!���Q��Lu]�2#�q�T��TJ�/� h0���ǳ�z1��=�+s`^Y�/��JC�/�f~�t2����[��޺�ӕ�D��Gx����d�30�e�*@4t�v~��n���>"kO����<t-��Q��)�TcP�G�
��Q`^��5��C6����H���L\�	���Ť��dq�$ݸcLV�����.�Sn�(��HN�2NpN����W ˟����^�qp���Dp�H��H�n�o���F�神Tv:&���p��Y��32��Ru��ʋ�x����p�o��#�`Ni���*� `>xʨ4�]U�xJ�AM�k�Ye��F�;%��`=�J��=��C�Ϋ{(haQ2D��Ca3�XK?cϜ>0*U:��{��y�Ц�;��44	�~�]>���,��M�WtMy���*s�,B�lJ�>��:?�ֹԖv�.{�����i7T��M��wcT�2m%`���3�by�#9��O��a�ԓ��G�Ї��$nB�� �+]jϔ=ꈐ먚j��-�^ihb�{��5T*�$u�Ǟ������窢�k��`r.�)m9�)ʽ�&K&܇�Y����/ ѧ�Ϥ"{��T��&@4�Wݐ[�.��xsVP!����'�"���0^:E[y��Y崟�������U�q���l�=z�0����Jx�i�`9>ױ��<��K������JP]���s�4��|p�D3�{s�L��dS5C�p����R�u����@${�-_)y������$�3�D=���s`�f��F�KB= \lm�^b&�b����幏lJ��|��לc��>h3�4�lg?|@�� ��Ys�A6��B]�/
T'*��$��G��&2��|EޗM!ݾ����19
T�K:�=/}��� &2�s����HY`��0��m����xF>���'�-��I�n��Z��m�4��/!�����s�K�X4��^�	���nt�0������(��\Z$�H��8@��~yT���ON����7��2�����j ���Zn�!ɐ<��C��/�{?W����a?��nU�wҼJ꫼}jB�!77��Rd���ЇA�pv�xei�,Z��|��:��;ͳ�f�߇i��.��O��9qS�ј�=�k�w0�j`�m��a� a��@7Žx ����Qh����"�"H��R��ul�����֭r�j*ȇ$��y����Ƭ�:O;��ʫR���5g�jz��Nw�3�/��e���
Q��x`��ӠS\u}Ո�����4m�8�������)�z7�S���u�,�$}���.��%�d�~��*�MM�Q)�g�S��H����se9ϐ�f�d(����!���'^��^�Y4��7�h2h��D �Dv;f˂�f�h=[���8��|T�-���\���83GpӉ��Pi�^:�����u������`�?jh.�vz7�p���lAg�x�=�m��K�T�͘E�>�"�g����z�3+�2PCxj�.�a�!`#�@6'|pd���/b��e�`z�9��5��2������@��Fc�O	x/��"�
��U���$��X������zv��Kt�^*@6�$�Z���¡�`:?����hq+���/�EP����=-,�S	��L�h�k_XG�d(�j�!u�V����AI�4�h�������4����Z`6I�^�J+��pAҕX���&M�R_�
�8ky�,��Ԃ^S��r�m�{�K	Q%lv�l,�F��d�Lۯkg{����n�H�(QߞxFtͤ�����3��/h�*�=�{���dV�6���Q��N�O>P�< �H���#��%�V�o��+ńʣcH������m�_�)�9٤S���$�<3�-Tٵ}�=\4ε�r���D��tl���k� �)i��2�L|�#&2#@Տ'�i���")���!ӬY�KR�b�z�����]�ǛF��h�:r9�+e�����6� <f�G���t#oފi�0	��vc��j7��#�6��<�%��|ڔ���ub-���]�o���H��K�)h0�6�bF�r�٤��ѽ�6i��ܡ����O�O)}<�9��d�(�Zmjϳ��&ȣ���@5�!HB��5a>��Y��҄���R)5�#V�0'��])��|�����ha|�z�ߥ�Jk�2i7E���_���^��p1\�,;�Ip���Z����܂����}|n1.n�ä�堝�r  S.&ۚ��Wl���@�ׄs7�"#��cte���p�z�����vB��]�@dݠ�M��� ^�"BG��`Y��L�� ��|#��H�DV�L �e�pM2X֖�;�b��G	���I��$׼�8�@`�Y[1[�����b^ߔ��?��E���Q'��5���u[b�����ZsXW��=��LH�n�dVF�S�����?(5��=R�#�mH��3�Xy�YnZDN�Mt�-.߈���F�� ����ZlĆ3��&|�/������&�X����.C�6��Ņ��E�=B_��'kQ��	�3З(žO��ҋ>d���P��"�(������h/�4k��O�SJ��f�f٥�NK�_��$�nJ7���/DJD��Q��ŷ�ɯ ��o�sI{��M�&4�5G���g��}�q�Ӝ$�i�i"<�~ �fR&����S�(�R�C����ĊQXH��V��Oɍܨ���tQ����cDs�]��"��K>��g��m��s���y:/@ם|�&!՗5˺����}���ǡܵ!s2�Q�)���j�`X�m�j�����3a7$c�Ք�����Y1�Ͱ�1����v@�[S��VZ�����
z@mKW�>��$�K�H�t�/
�����i�de�:4m�z�Egh��t���)�����;$-�;�JKE9i�E�^H��u��].y��]\�y�0���u����ڛZM��L�R��֡���V=�Kd�E���sV Z��,� �l,�^���~���-!Pc��]�.u��$i�b�.4i��?n�>��m<'^v4�)���B�ws�Z>4t�tˍQ�~ysa��c,A�",��"���I���>�+�Fa������P�	�_����A�&���O�,�-N},���4zR�-�'�Ѕ�Z>Ms��q�m0�;-l��_�ӕ����P]K=vEus5�