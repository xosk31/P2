XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Yf�J�m�k�Ҡ�
�o�ӍV�E�$���͟���\X�]���߂��d*�A�"�`�+�	:�X�$�F���STlg������|���)90;D*��{�c��"	Ӥ�����궡�����+tĦi���Y!��1T������3��u��`�ޘ�n�k<$z���{���M�����c��~�S7�h2%�z���#g�A ��w�Q����%��1�Z�pQ��aԙ;*��7�Fy2�����Y�Z^S �����D�L7��%nh�U����ȃI�?L��6��^�r>�$JV�z��7ڿӶ%4c�����/ؗ�����I���P��! �pFM����kaE�S�M�#������� ����J<���۩�.��X�����j$p�DWS�zC�T��8s�G��� aB�V����7��w�ȏ#�ә3�b����8��}����ؤ�
_*�N�������	�S�6��: _��Jy��6�����*�;��E,8|+��EQ�m4'Zi��O�l靳���_�eXPq�!��6us�*t#qg��u�\KݯD��15�Zͫ�O��j�^.�|Jn�a�?�5t���˿��-p^�'�U��Ι5]��)�?���U2�#������	9�^S�p�Cktn�P�҉akzj{z�.݂���W.s�rL��M[GF�vIL�@�$�΢��H%�h���� ��'b�����v�r��-��
�W�k�:_�md�׳�g�Rkq&ކ[v:�lȚXlxVHYEB    fa00    1d70e�¶�5�CB��ʑ�����[䤜��H_��쓆�!q~����e���o�*V�Q@��o�m����M�Q���gm���@O.�P/����@�C\@�g�)Ş���x5��7����0Nkg���U�Avr1�ҫx��(��4���i9ΓY�ΰ���<�1����Z��D�����Fx���xr�;�ho]��C��zX�,F�?%zxo�������9ֳ���&k�*:B^e#�8�m>^��qc�:5���N�N�8'�Y���������a�eE��T*ZbE^��-[>t��ݺ�L�;)�!�J#WzY�4��)�!$��)��Ɣ��1ؐ�!�m[нp��'��ӗ���ͅÄ��:r�{��,��.�9l=ЋM�MN7^5V?lf���u9M����[l��͑��ARh��YF?6wx>xa,�2��.�Ei]��:3�E��5p&0�A����}d����%Ź^������`�&@Ŭ/�
ͩ��$v��D��\�h�Y�j-�e��aX&���	J��(�eW�|-���YEj�~��E�L9�1C���+G?L���*X���������d{�1o�:pl�|w�`��c	ND�-:�k
d��4iו�i{k{	Fyt4k�h}!Z@?*T���8c�p�V�Т�U�:��g����Q}6t3_(�?+z�I�H�zVR޶�1�;4�|�%f1in'E�*m����]M9l�����|?�[�+��	6vv�����r��<���[�,�O
�@��fa`�)"oS��n���Wx��� /��Ek�?<j����ְ��VU���cgο��, ����j{G?{�o��y�h���v�J���_p�y|	������h~%�uO~Jm��fٺ����p�
T����Gw_�E�2�i�C���d�ܬ�"�z�Q���nOfr��p��G��Ńي�	q�2���CP�e��!`р�B;fDM�Xc˘��$4��:�k
~?��5���?�չ��a��G��c4�68�r�P�8�1�Pr����-��P�vx!1A�վ��)Rj+M6
�ձ��0�!K}�fI�խ��;�m�/�05�)��#	�k�٥���ίkx�vR۾n\����~PO���D�w�^#M��E�ЛV���sf�ܵ1V8W�)���_��^Zѐ����Έ?���5��b�/�b-�8���u�\7{���u�3��������m 6/8�}Q�y1d'�+J�>I�?�.�#���~����b�e���ݍ�����?ۆ��)h.�oF�!��h�G��T�Vj����qY
�"l��]���wa��3� =*��v�(yEK>�_s�x.�>"E5��E�.�v�EN�����������}/}JiQ5�#Ka���ĽMRVX=c�]J񱚀���NBoA�i|H�MM�����DMp�)����R��h@7�����޸/�U�n��2��$@���1g�%�����n���6��_]�S��5y��>���p�q_�y�����e�@��` �#�_�A 
�`%v- P�.&��hP'd}Q�>733��1ݒ���\�V,��S�t���g���LM w�Rҽ;��SP�����%�'5v����C6_�	�����X�h�m�]%���,������r�tM<�a1����]d௪MUAKϫ�xFr��K���o��.3.����\Hf�r����>�`��Ѱ�+0Ϊ����,�"Q{�2�r�8f��˭��� ��z���1��l���Q�ѐ�Q�����/�J�f�h��l������j{>x�H1�D<Q���qo�yO{-� w��C�/R�jB��4?~�y��]�7�4��o���
-�MZZ�I���U嵛❦d'���OҡD��U���(Y�24X��d�){���F��Dgqz�P��B�X`v:�0 yJ�P�[�\.�Z�N �;�2��_Ҩ�a��V@�s\5T���	��!��	��t��F"ޣ��#� D��X	��u������|"���Ë<���Iь�wկ�Ŗ%�g�ʪ�[UǯT�N���)�Y�<�R��}�*�U�;��'$VH*�֖�R1��
�&ӓ9�/��T�M�Wq�v]���Oc�� 	�a`��v]M|$Mei���O��}�m\�W���}y�8���W�,)i�[�'C^w��X��5w���@!��D�Ph��G�i���ޥ��nf��/� 	��6ND�ce���ɯ��_����u��([j�3�+M�}Q��H�m�~�`�&���6�@��v�+W-'������jʀ#07R��FI���F�@��1Ӹ���k�<T:+��J�[�n��(���E��X��~M�h&Y����NCj�����0��Pnz���B}�'��W�7⁨��I�&���\3L̡2���,F�]�X���M
")=�-G�]s�c�^�:b���<p�S���ݲ��g����٬�`���U��S�Or͠���}+��Μ��p�����(TOc�N��!<�*c�ݐ���=���z8�hcu�|�U	���!P?~|4�r_��c!_O�IL.jK�U+�U��Z��Wq��[���z�����*5lD*Ժ�i�8��t6�˦�Pn:C_���� �����y�d�y*��!ݨ8����$G�F�0��I���Y�3�~9(�%Rlv�/��.# �}�P�w�i��2���$�����7����7��=�0L���1��}�]J9EZr�i�>e��Z*!�3�4Կ���0�f)\㨈ْ�G�Y����iF�X����t5g�Ң]����/`S"�!�ߩWw8���=cT�dKW�rF����hC+���c�lQ�aG�fE���x��?x�!��eM�\�u���%�7�V�F�x����2�PC"��mg�jM�.�z�*s�cwI���מTd>�ܷ(�Y�ҧ��V�~��Mȏ�����5LH�v�UL�Sq!
؍ �R_=?�����zo�)��ތ��3l9��@��c_��88����2�&|+�A���Y���Sq$��EL��iS!<�t���ە����G�8����এ�2��+����)`�(�K�9YS�s��t��<�z#7�Y����zݴQ�o"G��%�dӏs�������b�gz���3�M��x4Ɔ2u�q�6���c��6_߷2�y�^9���������,�Op�=����9��Gcw�s�2�*��=���ӂ:�-[B����1]�Cޖ�K�U�����p��Dn� ��b�[xxHf��x��l�����n+�`��i~1<�X<g���e�ҍ�%ߘ�E�B��0T��k��xF�1�V����������ȑ|��X�4d��i�վ�7�=���>���}�Q�x��_#���Io�	Ù�0���/� �B.�0�z�'Ѕt_]��ׄei{�� ��7o�ia81�.�l%��|^�������ҳ[%8�w�7�����r8υ�G�B�x ]�"h/YS�E���+PȈ7!|H.Qi��!�h�2 �k6Ը�K�^���r��D���
+�a�E�=�PА}�`B���&�f�a/�ǌN8ʎ���B*��hy�si�� �����s*_U{*���"G1ktC^ �d�����p��C]4C�p�E�&��̕Τ�t�O��56�x2��8,nRL?C�Ƿ�w6�r�!�o����u)	�����<**̦��b��B�F���-�Hf҉�w��1�dr�]Y9@4�BI�7Uf�:��b�iJ��Ԓ��Y\�n�}��.�ڲ}xz�a����Y�]�L��R����%]�x�A����fD�?�=ѫ	������^�����D��]�Za,q�7��\X��ϳ���8LHQ�K=����*�>]S�e����1_��kq���7>;�g��7�*�s��ĂB�a�a��@�z����1�xɶB����V[���gk������@�U8v�E �"��DO	������1q�	"����˅�c�n�{��1[����?P��%��x,���j�l����۠�tf���]�m���u��G�P�;�A�jq�ZO�)��z7� �+r ���Gt��ӻ��7�E\�Y7Ѕ�9��C����A���}�7��Z���� ���;>�B%���)��'7��b,p��$2RwC/��so!�F�cD~�ڝ=�(D�#2i&�x����L�K��� 7�i��L5���N��H'�Nw },ͧ@�y�)91�lr	�6�
=�v��7�:_:~g�י.pF4�x��������sIl�L��D�"�_A`]L��!��z�h�z&bI�&;h��@b�h<R�eiO�D�����>ȞP�/Z�ZYv�cW]��3+bS��sSоtr��=�P�V�EB��.���or�������(+�d����I�78���0���ً��5*Bn��ua�ݟ9�x��j�z���Ȇ��)D�S���g�s��p0�E�B������,w��̒��kM�Fօ��0���>N�>V�|���!XԶW���	�!Gx�пye�C1��GK�K=u�.�j�5��n�qP��!�@�n�
�#���	�Aj9�� �s`M�����
��P����R
����$�x��P�;cxR�[o�!�Q��B�:*��[��
��Bn;_w@Ʈ���P��`����(n����K��?8g��U��L����>ÈaI��%ʥ�v�!��+A�A����&aѿ�ƿ矪����H>Y�,���moэSR�q�� ����V��<<�?�hR7_���r咔��Am�
��goT;��ݟ�V�+9s.�9�*+l�A�I#i�ɿmV
J�p�A����7����}���C���ǯx�V0C�g
s��п�r��;�^� K>@�$���Pҭ&�K��CS��PF�Y�=ok��|~�c/�x�Gx���RM��k��#"�`@��+���w�=�ò�C�c3F@[3;)������W�}l��n{�p~ 
��ϔ�d+z1*�E�i^�1I'6�%���|G��|�X�1��?�.5ȋ��~��!�A���ͯ���%}�Tq�^WU�񡡻t���_m�<�w�Rv��]�8�U]5�`����'2���a���S�=~������V�nPI['�6[>I���6֥_~pw��q:�)�?'����\*����63\���Q vڔF�s(��Z�A*.y^l�>swr��K��pZ�c�5���=��
���r��̑bɚ����z�U�lA|Dܗ|��Ҥ*Ҵfqﹻ��R6��@�2ɤ�+4f����Q?~��1q�`�i��
h;#��<;	�̆��yG�n����\�-�j��Y�)���ͼtِTe��I	g/M<v��o���h܀�S��� ,�±�#�@����R
a�G��\��rf�~n(2����Q1]�ǡ��rJ{���<��hU5G�4�<u���$f���s� �~����H��ț�&�H�?C�4�#xG��(�<�M�8���%�)Cҵo��?�]�Ҝ�}�e"d�#��׋$ "�J `^�CR����,�#�(^F�6Ib�D��m�)�P>�)}$���_:���+qRt��wB��-��<��2�F$��{=p�򡡧NZ�'���U����c�l0��6f�����G�����X�B�? {�Db����i��)�p��w�-"��$�Du�߼g�<b1%Ѩ�KЛ�h7z� R�Ow7Y`�����#:T������h����b+�|�jB��*�3b��Q���#��&j��mM��|K��X|�r�.q�o�y��� îo]8�����(H�/�m+�LPg-U��	>D�~�y�cl*R�|�{�9�$T{A:G	���4��B� ��̽�4]j�CE�zEH��|�m+%`@�Tf*���&�z
�M:�{7Jk���u��s����G�ba����2__�"cI���~;����#��Av���D�����D��m73�_��Y���P���� �
�z�0�]��LcȔ�2�,N�s��y�<���������h����z,�yk{$oW]x�nc�9�ۚ��*��B>,�ZȝT<�|�:��aj��;�	�;����@,SkI�yDݦq�����=�gh�*#���:�0���]-m����syU!���ʝ�a��t������7������'r�	�:�%d�7�}�¦��Z�5<+p�G�:<��Q/Xqw@�=E�x%sf%�M�_�ʋ��j$��܁�[+TN����R�jƚ�)����A�?�}�[-h�#ǨA��M��*��6���R��Վ�#Eت�/1�@�o�o�Qb���aӠ�6�~l]9;�"w�Y�vN��*l��:�n��'���1=$���@�-H��̮3�8
�2[�y���P��ӻ����å�i|�T���u���uA�Ѵ�������r�W���g���h���'��1� ԯ0����)DA�A^L�܁�5UV�U2jka��I�az�|*�3ܣ�=��p��g�؊ر.@L�5	��5B���G�����Ơ���dѮ_�D4;$FRE{.Hܾ��D%u��D�r(��mV���+[<��H��3�>�f�1Y�H#�m�)�5��҅Ɍ�fY�8�M�v���>�S~��b��x�ۅb�1�Q�N�8K�ANg�oӠߙ��>��%FvS�bR������D9w^����H�^:��]|��1U��]���I��8"����2u3M�N�5�&r���̒^#��+��e�N�x�4݀��$W&���Kg�#�4�XV��o_���T�J�5�^]0�;d#e���O_;�p��ou.%�����y���񄂒��u���{/��e�kTn\EeF�̈́ؽ/��*R6�e5c�Nb�v�|�؊K�X��SoH�2��Ǉ�-[�`Ǆ~��LaDD�z���C\�V0��&���g�h���W^9y�$2�_��O�V�X�/�|q|Q�i�4څ�0�W�6���.P'�ҭ#D����C�֔�oV���a�-�zr.u�2$����<3Sv�M1�����5���(F_�����/LSH>/�fa'X���n�ud@��[j9�R�n"�����Sv.��ƞK�I�M��8p�K6������[��,n)2�7=3�WH?��Y�L�,�/��c��-RC�j��-{���%��D@W��ߋ���O�!��w0���C(�c�ɹ��'��$u�D��l�/��%�WD�q[��ez���j��.Yݩ�yC��*a�e��U�`���8io�,�Y����e�~R��DXdC��� t�k�?��#>�X\���\<"��͢ )�nZ��YG��������|�N�+�f�1�9���:u�^�@�U`ӡ�xԎ:8�m)	0Ǵ�4���j��tV]ݜ���ϯa�R	��;����XlxVHYEB    236d     6c0J���yE._-��p�	�(���Yf��_t��(/�ټh�b(4�\��O���wÒZ�����A���Ķy���4W��e4 z��)�`.�xq ������ �C&���%��k1a�m���hg�~�ن:����?��z�<8��i׌G�Q�=@��+ 1�5�C&��Y�-1(0�eGC�=��d�q�X�#t����;����$;`��dI�VN5�^�K�ҥ8��kU`+�,)�A1k�_�Y��/ܶS�1D�F�&9���E*Sk~��`�����)����(v1�����t��t�#wZذ�c��\)[��Qd�Šc����%fT��j�:T6�� ?��4�qę��`$�%���#��e�q~��/���f�v[�C�ȧf0g���h��.�j�k�ߡ,���@�Noj�0�YWN���C@�ـ�`�"�bC16R�c�<"ؚ\I�Q�i�[����G���?�)ĺ9�>���Zl;��V�g�>#OO^g��Yu�����OAN&hM	��:�U��#�"���)E�l�܈��*��]�Ц��4I�~�\�)�~k
'2l�\S�_��c�y���zCy�;�;��K ��CG�oC}gJ����\�l�+3����h ��v�Nذ�/&s�Z�W�'�p�1��1R�*)r�r�̙j'�,a�qyt�Wl_Fԟ���Ę��iy�e�c�M�M!����C����/����5-����,X���(�ȇ<W��ϼ�r�ɒ_;h����o�=�n��bZF~@�%�lv:tHTg�@<�\8���;���sA�y�CJ���)�`�q{�6���?�����F���,���ΦK���"D��JகW�u�M�0�Dc�B���I��4%��o�X�ci%+���T,\�M噐��#���ُ��n�����5��0��x������T��J�i
	y)��')��V~�¬��V���!��T���z���+���ы��|?i��:����r��Qc�vd'�m�gׁXKz�jOR�a��,^(X7pA)��6�AR8����뢨gU����ŭ�>�TMR����v�"^�4d_�I��%��P��݁�fg�B���)��)�w8y��) �n0=�[�q[��0�jC���R�
�y�J���r�HH�w��������p6��G��_DȀ�5<Fz��+�e7�О	�J���M�~u��(ߣ�X �HՊ���h0����(����t,�O���ځEIq�q~a�8~��vc=E��cRoQmn�vOG�q��e�g�X���/s��:T��#��jl�٨�A��w_~���<U,"U���3�Q�a�J m�7+��p����
���ʪz�U�C���8y�5M��Ø���HtH���tv�Aq� ����po�oD1��%f�p_!��\�E�ͣ�ۤ�����l,�E	��^�D�E�N��8N���D�,��+�X@eE�	��n|s����޷K�f����K�b�����0�mi�:�[ś�'����������-ܢxd�Fu^���b�*k����bI"~c�S&Ud�ó���B0p�%�,K*q�/��w��y��8`�)�?�7؂-�Jݧ_?�6j-cٺOw���8���H�F�{���7���;_�d���̲�l��9�X�O�]��!=�*�.ǊsL����~��a@���E�8�?;&�C�[�