XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��p�����a#��_�{���)�TN�ASJ�{0�(�S�1�8�����0-�d��53�dj\i��b�,��'b�����q�$�=%�m��$� eB�p#C��� {�'�ЍnM����Y.Y����8BJ�ĺBm����@���K˿H���Ȍl���tq	/\�D�,e93�Օ����v�dl�ZG��,z$���Ε��;�ͰT��*��o�%��rd,�pB�BH�j��1�N>���e>6.��O��?��O���n�N��ʤ#�~�B�i�!�L����#���2��O!�I�jl���;C�7�ُ�����n�8�`l'�_|��@A|�*_�m�um�,�{��Th��3<�ү� T����,�ݥ��U�c�v�=v~肀8�y��� ��MN\"����,�p���ty�i����{�p�v��17��CY�!di��a5]9�[�VA5���!&4�՞��F��V�>z����p�W H��QeY)����Y��DfZ-�OW�ۦ��~��*#W\����v ���.�q��_�{�,��p�9If�`���/���O;Ϡi��R ��p��>�������4�l��Uę�B���Zm�H��4���=�|��v�r�!��>�un
�]$O��~G�{c��u�}��P.�S�z5��:��=���D��ԏ
�y�.7:�h��KI!n�:)q�Y��Ǌ'��4���.DO��@�l׍�mf�}d�s_��M�����s�Xt*&���a�XlxVHYEB    ea93    1880{:�g��(��6�y3��v�l�Vj���ᓈ�@�5��%f����e}�>�O�3�0�	`�UoAD����wf��k��M?~i��t�%Re�kAQHZՒߡX;�k�#�}ޤ�L`��oP��ٸ�ie���O��k�s��W�v���bL�"v?2�Ħ9n��NYv��D��	jx=���T`}4r_1���b��:�ʃsqe��Z�����%���A&��Ww<u���`y2��ioarMF���<�%t�S��/�H��|������t��Q�f�p�J���%��r�e���.A��D{r���s쓎���[�Db��T����a�>�.�?�Cx��l�ʰ��.�H��Ύc_ǒI��g�<�6�n��(P�ħ�R-��j��?� ��3*�4X�0�� P�c�'�?ZK����Q��)k���m�pi����c�Y�Hk]��#��-��c�̄(��/ڊ�L3
ٟa�m�Z�n]��B-��(-Q�IOT�G@]L����8Vhݺ߰|W��_�y�����G��(i��Z����*���:`<��ʐ�w��Bd_���0ʖ�o��t����?P�82���\�e�ߗ�!�3(~ف�[�s�~J@�Bs��s\���C袾zV&���NA`�5����{jU@���u]�B%zS0��@�k��s��,��b>���h�e����c�h}�T�>�o�a@�i�'at�uc��~��1�԰C w 2�E�ٙvCT��u��=񰀻�B�><��Sr����\���cS�^�QNu���'����6��"Q�W��*D��/�Q�(�Fb������⭔��O�K�y��4z},T2o:O�!7M1O����f�$rj���+%Wz-��עe�`���{A]'�-�?pX��8���
*V����.ld.�!��^ۊul�^i`IO�8W�()p�*�3�I�c���2��K��Du^�pS�R��������E(��>���C�o3h�����W:(�h�<q��M��^�PB��<:���xO�3�TM�B`$e�=yQ�����Z.��&~͈WPf-^�4�<�Sr�����t(pd�ﱬYrM�9�r4��l|�J%�-:�F""ӣ+Wi��[_H_� y1����e�]թ��Kn%j�ӿ�3���k�P��D;{�F��y�h��,�5�9�Ƒ*��=�VwJZߘ�,Z�H|���E�_��?�6-f�B�L6j�F:�꒎~c�p�.��`�}��5~O��~l��C����++4󣻔��I�{_sra�H�"Ȧ�L���/��y��Qۢ��9�FT��q�%[7qбW� �͚$�HsG���p���tut�	e�;�粨"��ɘ%x3��2F�L�?�a�e�����7��@w�W���b�����b���qI��g����gt8�=���4��oQ:��QG���=ɭ9?�/a^g!�����(\b��u�{'U�ۤ��w�EI�����8��J׎�ݴ��X�Lg�h�$De��Ro3�λ�0��b{J�����8^{�j��3�\��c)k�����$e2jH�~�qA�؜s�Z�
C��F�#��q9}�%C��!��9�?a{�z	q����&d��OF�FS��5�4$M�l�W�B9C�Ҵ���V�}aj�"�a@h&���T?.a��ŵzC��Ak&����r�-�V�7�P"��$��7�
,�i��Oo�ⷺ	jo��jlFx��zx�T/=��M��k�L��ژ�K���N����J�w_k��|����T�)�X�Vğe��"�dQ+E��֒4"5��8�-l����c�J(�֟T�ߘ#�]��:�W`aȨl�#-Mmq�gh]�z�-��֯��\T�:g��� �� �D|�ز�:�K�Z?M@��v+Q�W1�[��m)Ĭm�E���F���7ۘɞڌ�j�nTt:�������[�E��:��zK���b�e��^U�*�JY��/��P18pp���,t���,q�2�����H��G0���g��f�/Z'�B�*|i�?['�x�f�+���o��#��,W�^�i �"�۔�eTt |E�*�������)�%�ȵ��2`;����j�00��%�9�5�0H&��F$C:���e�>���̪�J 5YgytP5�~R������Jps�)+" ��fΈ:
��h��,���9�g��dG���p�o[ƝI�V�A:ƻǐ�:���0?�I�����2�v16E���ۻ7lK��J��++6?��{�ū��9���`'ѡ��7���DBaD��[��l4`؆�r/��ZyXk�*l�x ���$5�:}jT���[�x��l����1���M߽?�q����gF�0�9��ص���a���7��d����e�g��\^����+���t��
?�e��v�틃H����'Ʃu͎%c{�CV7A���C'��)P�b�?�>�zb�F�\�����4gq��EJҵf@l�%&��t7����_o��3gӹ"ͧ���yTD�>��b���}F(7�a��U�Vfe���k���$���wU���tyi�m�G\�O��Fn_������e������zP��r}�Y?Ǖ��r���D��bT�;/���)7�w�!<F�{f�!@��*��!���N�j�J���7?xn_�$Z���?�az�̈́�j���z�wAH�F԰.�O`��C �3I�A��6^KC��lE��N+���C�<����,��4Ѳ����q�2��<�|�T
��"	��Eڗ�Cu%��qj�|d���)�@P��j���Ҧ�8F���8���g�����O_Sc$E��M@�����!�0��P����y;i�
gO�"������j>Oc�CX�����s�����nx�������%�Z	�ŝMJ�rxJ��
f�H@��}�5ɝ[�\Q]�����M�5���#5 s^>�bnZ�a���CG4�]Y��gX7YR5�J��ڎ��utyWY��g�O�M���sl�M��
k' �b��v�^������4(��(x�R�+/N����d
&L�}���1��	��\��  Aa}+�X˓��o(�l��P��!�>D)Q�cĦ�`f{~RO[h����@J.�	��z%(1�I)~Qv��3L-�F�
�e+ܳ�{)gT%�����i~��&c8��#޽�:ϙ0�	��$�q>>T�A�f�,1��؟EZ���gGQ������/{ѯ���"�J��4���Q��.;��m��BG*�����n�
0]�D���3���(���R�Xh�Ѷ"���]���1� xⰲ":i�t�PTW��po�w�\"�jLK����;{�$ۘ�T�zE4����ip݃��P����~qMpߢ���a:]�g�Q�i:���3N�PfH�w/_Wp1��-^��~z�Ϧ�G�}0_T��'�;��Â�b�(׎L<�1��5e��}��C�V��x͹�'6#\:���1@�W�*QXd�Bֈ�OX��Լ�eW�5��T'Z�Z�H�֠�zy<��X��6��/��7���>��<6�?��~3��c��&��1_� ?ᷔ 6�V���Y�O>WX0�����Pc<kw�"J��O�2h+� �h?�?PJ�E2,H�5b�^�Y�en�!_�������g�U�*��ZE�A�n��P�\G����ʮ*�z� K�=6�upw9TTJK��t51�0�M�8vQ5r,�5CܗBB&��g[CU�s+��3�BC��g��Y�r��+ Ӎ�+��d�#w��=SX^s��p�eh��Z�JQ/o�{ͷ����ȇ�L��{�WEX�P�*�P:q��&��F	�f3�<�D)�^���^Z(�o�R�m<S��[� ���9.ߌ`+w{�!�D��ql�}��aG�jE��E��}v���TG�F{����� ~�?>b����Ůi�N�B�?�BsӦ��ez�p����D��ߎ�5q���qR,�N�c;�|Q�d�F��?j^�C]�,2�\��`��!PH�Py8.4B��aH�M��oD���ۀ�m�^3�E��yM��>����,���$0##s9il���:��[;���.��
` \�J����K��cNf}lb��Y ߣn�������]�
t��9��{���]^4�����k������$���pO�
м{�U�Y�յT��j��w��x��z��m0�}�Kn�Kp�� ��a�P&����!�\�V~�L� էJ�7iM������0&ѐHo��Fɴz��_h.�$o�T��r��'����;c�
�{z%E�z��_��Rt���n�3�����N9�?�K�}&ٹAn�r-3��n���y�m@��E�0 ǳ�������K��'�r�8y<(��;e� �pl�&?������s�X�H8%�"��O�sGn�a�E +�[{Qh?�[�y�{��>�"p�X��'��&����� y[��G��-�;P�T�P�el�f�=0L(n/��$�~����z��Q��;}�ɦ��,v��m(�����+�c���b�U�D�)H��m{H�g�-!����j,#�p�
"��Ld���v+E�'�Ov��3�nLjx�aȚ?��\�W�������tvg׭2	�s�Q�&��ؐ��%eLvQ�ku��u��d6߂(�څ
��(���~I�s��t��f�^�z񹌇�^��H�OaG����=?<��E�Ǣ�Xȟ�����R�[�|��H�?�|Mק�A@���r((��c+X&hzd�x`]tu����?o��-� S�9�{i~�H�T #0�3+g#3�6o���(ֿ�����@�?X�x˞}���'OH��L��|�Nj�EK)��;ހ��l�G'Z�f�/��Y�x!#V�şB����a��Q�Y$�bI�NW�})���*P����nsZ~�ei��
x�
Wb2��5�;���vl<��pCBY�N�Q=��%��X����W~�{���Tի3�������˱��5�3|���T_
xޞ���GQ-'���nȖ{�){5�BC��x: i�<0�f����z�#Y]������>��=X�VP��\_�⒢��}��&X�
���w��ƴO�\��G��րbN*��]���}J8��8�蟟� -����^�,�-�ɉ�m�fz�ɖ�� ��gXd�����3<S9Z�L���.X��5�����H�U����Y��ߟ|�Ư��U4��h�qJ�3�U���O�V�-���c0�h�������sF�8TfU�9҄F�	���R50 Q��Ķ@�
��{�"V7�n��h�NM��c&�}���&�L��V���T��ԱI�>��ݓQF%�Np����2Ʀ���=;?��+r�~;[�{(�Guʎ�Z�d����4�>L��'�7Dw��>�AF�S+��
�^1$B��j}9���W�?����][�ߎΠVZ�N��魊��ٗ�c�!ԃ@��<!2@��P0w�!Ej��)����do�cV=\�.ron�sH��uk�!���i��a�(!�t�-@"u��t��D{�m�[�{;�-@�_կ�3� t =;;[[�W���B�bé�ċ.��8��o�s'�<�x�w�$����#@ٱ�?��|�����B��S���,5b;s>�o��b���gX�v�ٽr�ψ7�i�w�DY#�æz��^�F&Ք����p��s���J�:�^.�g$i&��-B�K���.�:����mD�����F6w�c��E� �_n����G�����{:��J��l�UA㔠FG�KL�@6-E"u�x*���U,�̕�9�}v���ܹ�)ԋ/��s`]���=�� �y�f
�GB�ͨw�2���մp$]g��d[>WWB��.��E�,��&�Y�K�~��&i8�����.��<S��(U-���!b�!�P�uq�w��X���$rqoDPb����`J�pO�x6��K�� �]�7}^�*�+���E;.|kR.%�ڈ)��Cgg�(%=�	�7�b�P7B����_t:ʄ<�]#��*=E��Bjm�D/e��SY�O'�����jզ �}����W�nt�&އ����ҷ ��P�Sr�[� }$��o�)�h&�����a �n��e��zAR���v.�O%�K40�4�k�?HX�-�d�.�ID�6Nʵ*C�k�^�(�ё��mG�v�|�	���!���2��D��~�+{�˞M)'�����w"Z����