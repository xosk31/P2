XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��]酻�U.Q�V	�O�ޅ�ިj���ꄭsr�ܽ�,5T`����u�����&re��X��;k(�"jXi�e��d���<n�;�'�57�;U�B�!��t](�2��aKY��M��zF�*�y䯂��Z�%Ņ5���;eii,Qy3�ؙ � �d�xCaIc\���	i��G�qW-�.rn�^=��[�M�f�FS�=�ϒ�K�*+ ���d�*�V#c!��L�f
���`F.Bɔm�zr��h��m��jn����X��uNoX$\BPLƌ�����{_=\:WZ����O�R�v<	m��%��/�P�����5_���:g���i�:��HI}H� �)A�;��L�z��MD�Rr~�n�Bl<Yx<]��R�> �n�Ǥo��bGA9�e��A��R��2h��CK+��ų[k�õ�:��,í������W8���H]�KW���0�<�����*�/�j��PQϼm3A�NЭ���	����E�.���f�A)�?��[YS86.���}ڗH�O�!X����ԧ\�/����B7�>Z%!������G��|*�+D�k�t&T�i
O���\��I�3F�� K6�l�i
�4x��HP��r��
"��V��	k�Jo�]j������j����؈�_�ż+��10GUu�*�#��Tn�w9S��r� �������v�(��p�G��>LDS.�f�F9eH��u��h����K����U-����G��^~��F��f�ݳLC�y>H�X�Z��^�XlxVHYEB    8388    1740$����r06��,�����	 ��7��A���'�d�Y�h�$[ϲ/�;N�[�w)��+�y >���zgf�5�}w4���t�6m�����\��7�Ck����$&�P�Q���\�2��-v�����:��k_8���?`��2��"�X�>0�l����sv�7p>�_o�#E��=M+�7�*�e�{zY����%�z�c>�;W,�0�����(��\��P�;�Ij) ���o@��:��M��7�	�����F����ʟ��a���,&W�@���(�HoB�[/�*ȡ�55���xo���?A��|x�ɛ�q��A��}1O��-U���m�䫲��_��.+�93X��#b�8���q�.��EC\y�.�fᘗ�  (�U�s�ց�ݺƥ
&bu#�E��e����'E��+U��@7���c�rƠ!�>Dٍ2&}Fw�͝�O�Vʯ���O�R�k$n��\e����k3�B<ǦPrH��h��s���T5M��'��S�}t��!��p���݈os�Y�	�H�@���<��\�Ϋ#>�YviP�����2� g���{�!b�����)̓�L��mk����z�U�#o�,6]b�SbH#�t�)����v�VX��"��V��R��x���zI��-hR����w�yo7���1FZ}Af��Ԟ	Y�O��(<�<	h��4c3Up������3!c���T�RV�qz@���ހU3���v,4��<�fa�6����d���(��	�Z��1O0
w�Xk��zQ�I�����c��W�S�E
�_luA�n�`���֘��]��,m����!�*hX��54�?��^f�N�W�Wڠ�zg&�����/Q��E��DDU393�!-��ں�g�H�z�TiU�X�'�k2Ǹm�p;e�DB��*9�Z:}��)���"�4��l`��:S�&t��P�g	�ao,{` �[xv����'1(��_5t�b�4�"��O���ܾ6� �tc��~'{�Z���G�Ե\q0�N�xk�������������ӨIYǟ�ɉ�jK��͖ڎ�?��9ՙ����2S��h�|��p�K��y�m�I���bAę��'�����.{���U�ӭ�C���i��zB�j�~��#c$��ذ|��k�;i���� �1��:����c)5��`T��`rnik�y�G��.�W�9��"���d;�����һ+�Ft<�,��n��m�۶��(��x@�Y��4)��y٥�h���Qg�*�z��\��'����!L/o����;^0�s�����H�o��<'�֨�Q��C�]ّ:� 5��	�jq����8�x���w�-�9�*.�wQzN^K'N��9l�Yb���#�iE	g�-�{
U�R�Л�x�J�@���3 �-�3k��b���ҹ88H�2:B����;8�H�i���'Z;t�e��ԯ�<G�
1^�_�##�c� Z��(g����&��Y�|��̳��o���J���2�_�Y�3>*]���-�b�\c/l`@��TM�]�+���EoP�U��� =4S�������C	�����*�Hx5��O���)�V��b)j�Y0{
�ـO �]!��"���BMM� �
j�|Z\K`S7�\y�6�}����
����.�ł���h�&,d�v�y���C)�م�2X�ٓ�"{=��4�j{<\I�_�!;��C���X&1A��x��.�%����V���a����2r����+�W-6��>8���u���O��C�SD���w]�����$��=��R�4J���������Uף�-�n"�L(�%��z�I
�w�Z�Ɏe��C��^�1dW�޹�=���	i#��Ę.S.`��Sh�y==+�pDA
�/MIm8r�EB*w; �2�7u��nmm�o��+�D�6|޶�*�KMG���~�Lf*�fߟp�PL�9�y7�ܹ�>��X���_��yLh���_}�/{�8{���J(<6��$�Z�eVx���W��p������5%dc�1xA!�5,6�`����3G� �� ^uu)����m�g�d*?��F�~1��*y��N?����GLK�>�+C�\e�w�`��lǄӅ�+� � L��/@�� ;��9��Z�ö��"3n�7�^r��8���z��.��_p<sJk&�B*��r���<d�j������6�k�-���j�V�
�jwI����p!6'&��>IoY��S|��=������3�8�Mz�y�'J>_���WC��1�3M0-[sVX�<�W:0޻:�0�]���}�r�����@A���x�`�>���4�nGV&H6բa-5?�Q��CY���C[)zb)���vC������Ҹ��U�?���;��͏L� b�q&�Ձ��A���x-�Ე�2�{D!�W�=8J�Ϡ���
�7j��`8I��TyÖH��c��0Ԙ�.��
��z��NEo�=C�F6�����t�A\k�w�{?�d�VTP+sx��6�S����a�m��\�� �	��H�0O�����l�V5�����r��-�.ZA�Q��{��a�l:����c�	�W.�� S�CK��/+i�#S��0�p��@��|i_���drn2
�N^'����B�mC�Ҫ:!|"_eT���a�:��cV}�]͔)݋�aiUHm�����W#kTr�w�����d!Ϙ"K��O��J`=%�w��%������ރ	6���S��=�S�C�_o����<�Yg����Z'�͏����Z~��U���&5H�P��ӧN�@��^���Z��]l��q��&I���&��瘇�C��{NK�2h�j`1�՞�̘6�i�WԕW���50JmRݍ���s��p
@Gu�.xm�s4�xÃz�8����|&uX(u�~Q&��̙yA�Pg��Bͽ,��qw�@��˗p3�!���}M$������f=��/t��n]U]�i�1��S�ԅ���Y.]�nq}zM�����疉��l�iձ���<�fpȽ~b�-�nx���h�W?�4�T~�ҧ�n�����W�����˹��r�*�w���%���bN(����2�n��X+4߭��.�MWN�*�9T� |��
��!WZ��g�+�
�k4>W�6�"�R��χV�BE����.�̈:/��� �`�ty���R�lVW������w�h�h��)f�
;��<a��u�Ǝ�-�̭抪� �����h���KWO��X��3�Y����T$��ϧH+gT{_�Br��@1eQ�p����eE�r��2�����Q��������yX�^�b�$n�[e��o���D�@@Ĳ���������.��8N:i�/F(�7��h���s���Ft;e$����tE��ؒ�(M� �c��{.��T���PiC�z��c�����;����.r�	�����G �&���D�f�� �!�8hp�����c�S䝨��>̼�b�x^G���`T�v���E)D����F ��]0�E��d�(�g���0o�e e8�Ze.���KjO�jr��L�qAʲ�4�"[07�ь^ׯ��H�3!����o!��Ym&��(9[�c��#�1Ͳ� {]�x�5Z��d1y=BX�bRb��2h?��'B.H'KuS�
F;��
�8Ε���$����|���z$0�>����kK.,�LU�u�C8>�M��� �����!8_V��%r���RO������@`�֚��i�A��JB%�f,^��?�z�M�G VeT|QxEa[�>[�@��Ʀ'��
\��b[܎Ֆ2ꞇs�������?�l���/�1D;8������-#��K3���D�Z=ہ�โ����r8����P$���S��8�pv]͑����q%Z�>����yN��#�θ��̓8Rl=�$����T���%�!� �vM���P�Ke��ݵa�8hyS���΍��M ;���rSܳ�'��)W3}ة0�?���-ͽ�4�Ia��T��'T��ɗm��u�d�@���͔�B%���?}�-e�������s�?�`�h�۝��UPc�Q���AX��T���V�dO�!i0�ʓa��z�,�H���K�2��
���#���������[?呾ڮ����G/b���a9�h�'�%�!P$3<���%|Tcr�n�&�\�H-�4s��'4��b~e�Z >���zj��L�7�-������O�/�!%�9:A�������x8~_�ŏnS�0u�P�ڈ�s�ו�WR��B�h�kOB�M�4ï'�w�^����J�Ϳ��CצǉZ��֍��ĸr���Z��oVJ�+@�m���$$J2����l�����N��V�ZzϽB�.3e��IeQj��ý&J���+�|��Wp����y���N>:��J s���{:A�_Z��h*~�bKA! ���mC�LI�2S��\;↤/�����:��k��rr����|�"T�p�p﹃	f�ŘB�4Ѷ�F"w��e&:�F��!�& _U��YӔ�����^�c����i>�Y��2(�/ߥ��NṼq=�d���<����F�
=*0a����Z ��j9\�O�Ie@���E%��cf
;T�v�%1��2@���:�g��חB8�����'�c�"!�U�'{#���Ǖѧd�/f�R�q����n#���X���HFo������Ξ(ЗQ���A�V�ȃq�9 �s2����`����:ٶ�&yx+���}18��[�Bx�YUeC�!Ln��Xr��ɷo�hX� ��ٙ�"�,>�j�	��}��>�m�c!U�c2��;$Hǟ|��uWf�_�0�CY����� �r��5���<S��d�}��ek���V6���i�Z ���:>+z�)�8#�?;Ҟ �g0L�( S��!4�x�����e(�Z�������z�6��P�^�.d>�muIZln�<����,�$:��&�{`SY"L�0���Z�,
�RV8�o�t�3pA���R/��҆��˚�DbS	�7���i��3'�^Y��E�$�U
�j6��l�y�t=Ek3s���,���tT�N��'�[�D�$r����^�h7_�b^�ke�'��I��cBK� �$�V�.���d�|�X����fz��=O���e������FdJܦ�{O"�5p#��ޭ�u�F�1����]�hs�vP�����8G�q�k�l�֊�D�P���0Z��� [�N�s�ҦI�+p� 7d�(I$��O�Mj�m%����6|v���sZ8�/e+lt�ʔ��M*UϢ"���fd�$��%��$�}������x��������w󕝜�ǫA\:ok�o�3P�dPP�Lt��$�{.۴��;�������^�a��8z��n�\���h����6ED�HLJ0��5���>�z���O3O�܉3�����q��pP˛o\�����P�'u�^��L"r�� ����뼃�W�5���Q;TCܴ���H�h.�����3�a*u��da�\�|z�W�U���'n���3-j���ipLQ������/O����7�z������𑤹�בBWDc���n�������h5A�԰.�a��B�o��pd�}ۯ@�5�P!wt)���g6����J�؋��|�9Qow���`֯�_�VT�^����������a�_6�V�}��߸gU�_z{�5�,�V1���2��Ҭъ�w{3�@ҿ,���lT4	����Ek2|*!��� �6�>$s9&��z-�8��+n�ѺU�Vu74�!�����i�:~_Ͽ�	 5�v�M�^xCD�	32�t�!���2�I��]p��"�����ۉ�o