XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Ӕ�[+���[�S,ߊQ���Q"H"������kd�5~:���4y��-ZԬ��|ޛ/Rg�Π����p��ٴM5i֫�5A����u)���,�6.��>N�� �5������7���1[���撑�j de���U �������_�{�� �-�h:�D�?��k��`��!6�Hi?��-F��]*�#0;Z|������[��Ya�fd��XLZ:��+�n�ž�Ռ N�ZK;���Zh�Ij1�jNt����d����~�Fk.��*�m����O��7���H�Q!~���6I��%݅_����W��\�Q��:�f������̸�+�#s��@x����tO�/��ԝ�4-��Ǎ�=G���~;�6�Ќ:�p�K�<���^6C�"~��ؙV�ޜ�!���n�ת:���b]�V��r��,�S��ܜC�P��_e��qƸD���DH�40�?f��Z:^�|?�G��yje�~�r��?	�s��<0��y2[U���O�t���'&L~��R��b����*Uh�����Ȇܱ�Q�?`���&m��i9��ͱ.����^eQ��Z� +p?Qޫ[�D-I�(�����{��Y���r����L�3�vS~�y�S�NVh�f���F���d�9�f�#m��g�y��I�}�]�W�2ے��Nwr2���[��ā��Q�Ɔ�M �6��fd��sU3{I�qeb�����+�gش���%�)��U��q��w1�}Nu4�
��f����no�rCQ�\�O:D�/"�XlxVHYEB    1427     840i����Q\=��J�\��(n}�9��	���}R����mw��A���s}���{{[տ��"bOQ.�=�H�����5�giv��p���s^ҨH��M�<�����u����X�'{��ݚ�,6���b���/���%�ń�"/�|3��4|J�	��H���q|����a{%' Gu8�J����jU���VeT~����z��q7I��7q�hּP����"�d`}����37�bw�r����N�_���~�-:k�M��|�����*�k���?�_}����&����˝Gc�����"uI�w��W�wT�!�����(�PkO���x��uf�� ���wh�]���t��r+����<�=Ae2�E,���|��(���C.���;���<�|S�p��6ҹ|�q�U c$E�U�R�����q�iq�%�14�|:>
[��[��+_�`/N�Li�-뤇 u�� n[��1Bx���̡>�NQ��o��1ٕ_o{�q�@���ϟ����߇�صc�G`���MF��W��g�I�[�_��eL?կ��J���(�C$-E���h�ۢk�\!��i" ��)��o�X��١�d��M��C��g�nw7�p��7a�&Ӆ15��k�t�M�\ӵ!(�I��ȉ���ݖ����NA�6oV�ȝ1�w�bd<�7c^~�U���F5�u̧H�@��m�#�V��gco`�7�$j�)C?C����>�e�8�x�O�X��6	����^�]��V�P�3`VѶ-�%)֊y���^f���w�
<;2yAY�B������D:�p��!�h�J�E5g�6���3����UJ�VS���rU&ש֗!ԝK|؀u���u�
�Wo��%��O��VU�� �;x�����ם�R
�R�b�Ӝp�!0on�R=��b#�����oz�Qh��u_vy�ң�:H�R���.�U�X��r�����l���4�#@@E}�
����_��:r@�_��b�A���Q�y�*n����b,xV+��|9�V�~��f�[��9@`߈e���!�e�F� #�?�W�_�f���8������%Fƣy��O��Gʘ���%����&����D��2�}rG���bP����H�ً������b�ԋ9Ge����ӄ��� 	����ޝ�� ��u�� �ց���P��G+2@&KD��4��Re�"��i�}�Ř��f`*���&�:���MwG��7���UD Mz�Ǌ�1����:w���ƺ�mŒ��۫g�`�/�c}������<�G��xH��_��ފD�6�v�U�ԍǭ�ߝS�M�:�,K֤��^�i1�1E��G��3G(�$n��eϜ���[ѪAi����/�eQ�ޛCs�p�с���rc�J.EdqO��'Ux�.�ғ����ؕ��I���J,6��T{�!n���i�-+�V�
�9à-����S����TN�a�燜T�^��
�X�9�6���X�PJ��K�ý��}yJ���@��Cd ��J%Ӏ��:欖<���5�Ij՞a��^����F�ٛ�6�-�k][β��n���1�K<�����jL�y�wR�1�����X�<�gsHM���:h��� �$�J�w��o��=$
~;~d"J>wTt�����-8�'�S:HAS��>o�}�ѹ-�r��?h)R�_9$4[x��L�cP�cM�K��'�)CW[�����������Y��jOn9�\\���++����|�0v�L�J&���M�5�NN�����wGufZ����.��_uL�|�b�<�#�B��9F;��u k[(G��Tt�	V���k���t���3��,rg����c�_��HB��"�s�ݩd����6���h���B&ò'{}55�9�v/wg��='�g�5G&f��']S4���=�����I[�	1y�t=Cl�f��^�`��YRe�Sv�zq}� �XE�G�_��8������_��,ۦ4E\A95��]��K9|����6�ܫ��`'��h�`ZU�&�]�nA)�0�� �:)$�|ȧ(i��~a��