XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��+B��n�����6-�%�\����C��X�ed���d�$�!)A���ۑ�)��573�Lp���M��'�L�Ӧ�ff�Yh����d7s\�`B�N�������yК�=��׳,��> =F1_�.�J��ǹL��0s�X�����̾�k���0�J�'��^͌�؏R�6�GR���x������{H!���#@`h�s��K1��R��TiD���p�`��:�"��l�#�Pa�;���Q��CN��WƱ#AD#�N���,�ZֵVR z��M��}�*b�fI��(Y4�/�<KY~����(�<�?</�6��,:`��dLN�l�ߔO����!��>�}���i�}�O�����ڻв��OF�,}_�?���^�ݾ�ʩE�"�2�䄅�Il��O��JQ�k[�� �)�Y�g�
������� �S���)4!��r��w�g �sF�V%��a�?<SG8������j��(��{Ԛt/aTZN�t�Ѝ���&��yߋZz�?��FU')8�Jswd�s�au�9YT
��<&]�쪹���P�	VW��w��W];�#���G1c�ʗ({��Mʹ��A�1A�!��2u��"�(q�߈��� |;��W���!� ��D6`T����+ꠏX�h	yn�B|
�q�cc�a���m�*`-pk�1D!_od�*��#ޔ٪^�iMc�����-r��q�+;7��Y������S]dE�iٌ�D��I�S�LXlxVHYEB    aa31    1e40�a���ئ�yx
�j~|��u�a|��C����%H�/t�	�@T�1�z ��G�K��/f�2��O�s���(�(4�;��6;`,v�:�1!G'�1�:#(�7������Jl��R�'��h�]ڲ�ń6zoek�V�	�pG��)�.|i���oJK$&�
d�dӻ��|ԦY�qdp��U�f� �oC�#��Q~�w!�G!k�=0�����I�MZ�����I�f��}���G^6q�|�}��,�o�]5�y��eC�M��g����a�]�����f1����
n�6�<yF�P��\v��`S������r-o���'
K�M�pA�m�X
��|�.dس%���h��ze�ٺ����1H�-�.����I��Su����&g��	����p(4E������؇$���˕�!*2���o�\#8��CI��ľ�����Gd� 7�	��c@�hrw�.p��;.o�y6�%b��iZ|,`�T�e�Gm�9^��YυN� \�W��0��*ᠩ�;��bBǨ!nr4�Ϣ��f�̯{�ѿ�m�p\#�u0f��{�؜��`�j��a�/����N�j��q�IUJ���+�C,]��_)-����|yJ�)��T�d���Zn��>�b�6���}NPf5k��2.ɡ�i~�%�ȧ�J�v4?5Lzt�d��7������/Ӏ���R�{����e}�YU{���T�q}�s����ldb
Cc�i��S0rn_���둑Iǁ��=1��Y�e>�Xw*���1�F�$,3+�U�� ��s�4�,CJ�ThJ�����ڿvړ��%~Կ��>]����湳�z�����+�J��u���(��K�G������q~Dg}�r�k\mF%ٲ�3c������;.��6�����-�Tloq����9O2����-O>��)�3}�#q�p�P��qE�yiUj���ˏ9�tg����*�.5f����g��b�Saش��3+�-�6?�vT�;�ٖ9;$��\G���8m�,����[���4�|(h��N{�J�Lp��nϼ_�|jf+N]����2����É�HZE9� G��s��rƆ�)l/�;~��^�E�,�>:ƃ� ү3���w¬y,a���#@��,�/��Fx�` ��
��)1WJ��Y��(T����@�ƀo�۪���*K��07&����v�6~-]k4��87Q�)�vU��Voӱ;��T�֗:�,�k�:}*W�R�N	�O�[ʶ?���G�7��fdcH�o���0,��?��E�lC_ ��<���(k����R[ć%�V%s�s�s�qf���h<	�K�EK���(j,�љ�Q۬p ����jP�-��?���I�%��x:�
���y	�׮H���Pw����a
>㗡K����:*rXz�Α�	�8S�!m'\k�z_T.�_f��X6��B��+��(�����I`��L�״��F���v}
���c=��a�:)�ڽ��9 Do�u!�;�F
�)�?Q�9����#�=�{�1'�3�ܯ�v��O�-�N�F���Zq'Sԛf��%��rv,C�w��ϔ{��i��_?��Y.�=�W��l5�LPnN�@��p�q60�?����9��9m���NTo]�V'�����6h���p���eG*8y[C������ŕ��l�#4����(Op�.��t�+kZ���rYH�6H$��Ϝ��64w�.{�L��8�,.������`?�*򫻺# ��g�nf����(	�5�$Jqe����o��]l��x&BH�Uޖb10�mq�{l�۞�gw5�����b�qg��NL�����>U�u��y�����U�a �f��>w�T����K,��AW�WE��r;h嵨��:w����N����2dQ;I��������� 4�>�H���+*��������-�t��Մ;OĒEt�ȋ+gfi�I��r���Xu�w1B��������6��3��Wm���mw�/S�5���3@��r��?s�с�2ƛ����$���i��A�{��ȧrR���:���I]p?�zqU�hN�_�#.�{k��By�zZKF}QH,z�"���Ŵʓ'��ߠ����jFPA�-�o�,^����#/^��dE�+�ܺ��f���J�5��E�-��� ^)g�x'�6�d|�WZ�Ms���&꠴e��ʷ��1�-',f@!'���pv���2wtq�����#iؽt����1�.��QH�l&�������q����
�����НũSʷӉG�2o�uF�L��3�kK��N�cZ��.�0���{kͦ�͇$5ky�waރǪ�u��2S³W,I@o�O���m��Ҩ�8�X�ZoJ��@ ���lˎη�$*j8Hzx����~W��p�̈뤘R5h�6����Ԟ�F����6�e���s��Y&	���d�b� K��`]��rx=㨅�'��-!Ats��G::5ꫜ���.�beo�xsF�V����.��R<s�$"x���5!�ζ��ų�~(�5��瑐yӷm ��!�������J�y.[��6]?��:��z*��yXK�܉Sv�U�Y��W�ה�g�[Q�SP�\fc˝�z;}k���큔v��w0J���J�MN�oq�d!v��S� 	Y;Ӽ ��q$Il|���GU��0QXX�,H0\��^�e�F������a5'�>@���FXZ̬���L��1��(�œ��-mY��{�C�]�u�\A���f
������ l2q@x��I�1��j�̃��u&�Ro�>���F���DgP�9��n{���/���O��ݝ~��ӭ։���YJ�^�7�Wb���ǡ���9!��b8ڱ����$��j����
OJ3E�٤� M����G��]
�X]^�� �U�%|���^*~��D�(�VV="m#���k��2�D�#wo�[	l�v����\���R;�$1�S[49�k���5jCgiN�E���5�Eȸ���K�N
����F5�y!P���蚮{ɐ�j*���j��뫂�X����S?���)^)�/�&�̉�jv|m̈́A�ނB�m��h3�Cz���DW�EN+�/(qz���Կ�}��I�n
b==�l{�q碥��|Q�F�A�A|5Q#`vZ�,t�z�y��DNL;�'�
2�R���Ig�V��=����������?�@����@�톚Bq�:&���,�j5&E�/��D!�z���j�may��IL1�(����� ������y&~r�q�b|��#�u���l��jQ���ġy�c���N�j��@yi����OW-�2gϰu�wqR�Z|��e\I�Ff��xHݪZR&@.�z�n�V�X�G@��m�e1�����-U(���H}��IH;i����k{1]UԹ�}a��g��/�O@��W�������!*�G�K�?b��I��0Q�G\x�u��I�PP����!����G�y:8"�ZG4q��y����b]n:�'&�ѭ�
vJ�PON9{4��?���x{y�wi�f̂�����Psr� 0v?ʨ
��C���}�81��_���=�l�&�Z�O��2q���U뤛zr1�[�����N2f�)��-�P蕮���;��#8�RS���԰r��7���
�E��@%n�;�*
:+��!c��j�J_�1��U����B�.���ci�O�r���
��?̧������恞� ��PJ��� jZ*B0�U{F��"N��S�{��y6AK�%4d_���Ģ�ŕ@��-"w��U燆�A��b'{r9HFhѵN-ɼc�m?��<��pm]� /�O8��Ts�'6�,g�yo�A\��Mދ]��Í`�xS��GnP7N9�� ���
-di�dV�`��W�����44I6i.%��L5��� �a[G�k�V�������)h|�L�2�皞�2���?!���	����3-�mb����đ�sH�����5�yS�� G�(Y����I����M�2�-{��h�k�q���$\��S�
ܽ$֖�>v�9�[q#_Oz��Ck����Q��)�VV<hJ��4{(��=�$��,����8�`VC��H��w}Lسb"yx��D�����c�6��W���E�5��
K?���S���3��)���k���6:����4(8o��m�k����qß(����ˋ�\B��9gŞ�cB\�R�v���7�!P֢�#�ħ�V��խ�/���Iҹ�T
�j_	�A� �4��k<:�*�$9L\�@�ν�+.e$9�44��2�'#�C!e�sh�Fu�2"�-����h�9.��zc�C��B;ڡ*�u����ߟB(�2H�� �Pp�(��d��������ku\��	F�/���Վ/�M/�J�!�Hn��P$H������:嶽�D���$�"{�×�+�"�]�ӿalď�.4'�I����Cն�8}��&R������㰡V'E^���Ӏп\Xa������U�ŉU�-�Nb
<t=�gk\)R�HH%�����CqTݗ�I�z�F����,%����Y��sǌJ������o::+��\lY,�?���5�r������[�[Ɣ����~�b�B���'O�� ���j���(K�@�����C��~����V�/3�#!#�jnaW�T(o�bPlڀ��9e@��G-�i!�
��;c%��H��=h}������� ���<^U�|���;m�ǦW�#��_��
��Mq?� ?%w�� �	��J�8���[<�mS�NI_�/�>_0o�� ������Iӑk��:�R�9��lS}4��7�|HNN1埧+1����5�`u��j���@�(�,��))�ģ�z���S�����ùx�I�r��1p��|�@�E+
/��]�C��.�.ǻ��@냼ڢq1a��XK��1�~�I�z�߽������fBE��TN����@�+z?�xo���rr�(��n��B���V�w����ީ���Q�ԑEz��^޲�N�T$`�c$��yR%���y\�Ƣ��3}�2�0�quaM>h��'��σ5v?����uwI����툔�V[��<�(�J��ă��<��nq�lP2ª�^n��܋;��j��Oƥ��+-}���&G�0o��2���"�o[��Gr8(?�����@��v�_�z
����_�p>d�gY$\�?��)}(=�]v]@$=�Q�����VLa�+<#WD������b/ۭOM#�ԪG��+��&�8�g�t�T�����4�^{�O��c��(�n�L��pA�hv.���Hf�+'ie'?AL5k�|� h;�΁���0�}�0+_����N�o/'{����q���B����4;���ɇ��d`9����CX��9N�^�,�2��mq �Љ�0�{������%������<C�Qri�Hy��WS�*��٥N���L�:�-?` 0��vG�q7�=)`�h�;)\�GH	O��(��B.�Ft����iDY��?Fhx6�熊�+:佸&��Ȱ��i�M���RP�	��P��zܬ��A��`_W�*��a��y�_Pv�0��,j�_+�ޤ/��ǫ��	�j��l�8�"�.χۄ�ƵP~�u��
!�T�nǗjo�1Q�!lbo�̮IW����^�=�/a�?X��
 �I�=}�Gk�>F�gpS��h!�ڻ��E���y+g���`�L������� ٨��DΓLH�EQ_u�,���������5�E<5/5�Td<�]�\���#��*��~b��v���oT��W�ui���U���
<$zg<uʌ��MHwjN��\�1����0���Gk�s����R���S��ձow�~�7��zjd�8��ƾK�._���Ŕ��<=Z�X�-x���~I$�{$<��]/�X�&�l���q�z�0����-^ZP�/��Ƒ�˖݊�P��Q@f�cQn� �K���oD�&�'�Z	Ã�@-U��U� ��X�j[z�iۚ'=�d��b՘��1!���B�x8J��RT�d{�4�a��QwX㼹���<��V��1B��: �{��e��I��M��ÂLD��j
 e>\�c��=�NRw�ȗ�\�����GO���(o)����t�M�0�L�!_��&�)D��(T!�\a����:F��%13 �j�u���3p��D�J����\����H�ó��!1�+7s�R:(o��H��
C��72zmT���+�p]��Q`B��2��xZ���=�'9Ww� ]�
(�]x��i�_��M���E��F�)�v@�����lm =z�@f��X�SPۓ��=+(�I����H�AD0������A��~��c��{�!_�90�� �)��Y�ζH�v�	\�bg��h�-(H�@طƖ��#�A�?�����k���ctB�[k���?n�l����&b��Wּ��kPX�"�fS����V�R��3�8�B��$B�
�4�v��.��{���5]X�S+���3D����f�R"ڽV�� ��Ǡ�v~��~c5iO�Rq��&ؤ5�<�Rw�����[>([aCs߳4\þ�[�0�Wu���21o^X�l{C���h�O%:C�'�\K�{��3���=�YJ��^��l�L�f��v�h#��	�*���&���A}�:ǫ2"UL���*z@c�=MU�(�Nt"�TiMTF���l�	�C� �-�0Gm�Z��2�'�Y��2��w�)[BE��;RC�+��A�E/U��>i0��y(JX�o�s�P��i H�7h�ыCr"��ˑ2j��|��	o[xi0��[^T�J.*A�ڱ�8гrd�xpF?xO>^jv;�@;1�4^�]}ת�
GzU����w�us<3Xw Ӑf�U,�0��}��شH
�O�w��[
L�f����14vb�b�v���u��_yr��y9.�0��1:gr��J4�,�rhkD#���-�
H@��﹛Wq~�]p���Ƣ�4 �F�\���8a�Yu�9�"cq�i]?]ӵ�wCH6��t�(d�M��Ț#�);%ټͮ�1�sB�0vX !qd~F�Yf���x��"���|��ze����l�)��E��FX�m�w�D��1��� 1m��7�5W�xa&�L[�� ��;��|:��gY��\�nԻ�ݒX��E��Lt�v臦{�J*�9�������uδU\?�M�)��Y{ w.(�����GM��oZVt��6�l`�xU�jWG�}��,d�Sa#	N�^1��<Sb�3rL�Yҗb�f����Q�b2L��n6X4���b�X6)����5��XB�i���S�,7���֓X�;�����I"����_�dD�B����$X�<�A��c
{������z�79'�݁�;�L	f��f�xs��u=��À�E���}_W@�V
���T�]T�Ê*vIc/S�8�;>�//�.~���D6�V�$��9/��&͇�҇�ZG�1���[W�&WTx�!���%�Mk�X٠�a��X����D����+��H�