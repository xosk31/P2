XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����|�����k�l�1<���*^Sw��^�ƣ]'����ݽ�4��ۂ�����.���u�l)vEۣ�r�&yg^���12����1Z�����i֔-o'�������qu��*��bX����k#4|����ዄO�~�81Ȱ�쏞�9V1nޗɶ��R�E޻���;[��q:r��މ�Tų��-�������~C�	@��v!�O;a<�>������&F�&����f�c���5WQ:㐐s�N.?)����ϑqC��w�vt��T�0Ϫ�L�����$�H�#8~��C=��lֻ!�QS�?;�nE�����N7���qt.4Q3��[����O[���9��!�O1,��'�nѹ[b~-j8z2�kC鯂�GF��'��X@v���A��t�	uM����*nP���]�}����Q����f[�l9ד!�~�C����w?��l��V��ڏ;	�ӫ�*<R]Q7"����L	�[N(�v�;^���
#1+B��N����\�=���tČ�h���s�ZO�MNM�����`�B;����8���s?vt�v0= щ�m�M�S�$���� E	�ew��v`QF#k�^7�DD:5��^�Nǰ��.���gĂ|S��K��ʫ�?͸;ifv�X��������]�L�=��دe(�=?h���:篦�ؐ]��%%�i
` ;)�l�Τt��:�!lt���1����Z�B^�`R�)�$V�i4t�� $)k��n������XlxVHYEB    6534    1400�H�����S��=a�����3��|�\ˢ����������\��,;�i�������BFs����dϳT��z�AJ��QkU��{�z��2/N�!�CA�!z��y��_pY����AT��*�̓/n��r���1��xnZO~�]-cy��a�+'W�`��,��cr���j�F�-�@���J�i4ㅞ����]�m֏][�j��!a	�O_�tE&b�k�&�t���:���m���o���xa�hR"�xH��b�:�iL4T��K�`+'G�.��zcz�Ck�5
4������#�ǫ�b.9�u�=�Gs&?o�ȵ͛�t&��K����&W�B�q!�^�;�6����!��~��G��pb��<\,yA3ϒ�ZnH#����M�jV�`���Xj�Y7�Z��:Lȶ�1�A�oqV�'����Δ��:�݃_ t	U���;C�0�6RƬ���+[������D�ӄ���|r3�n���۞G�E-�(����B��s��QN�%����w���������*�l�\$K�v\q	��b
gq���>x)|����ɂ�I_�/���#��;�XȿR���RE�+L<��0�Oe�y�0�"}v. ��a��<��+٦<��p�D��[�)����.�=#��/r�_������c��r����ِ���D��X�P����S�0|C[��j����Z<'� 2�&�� ��$AH�7�8�.��aG)�b 	Wyʐ�-�l�s��!�6~���DB�1tY {P��h�bYγ?w������V��d�`��qJ˦�U�=�I�G��aQ���+�AZ�^Hmb�x���Ƌ�#�>�'{I%�/1#r�����RK����>��M\o$�B��9��=N-X?��y__��B��K��Vs��S��2"ݨ;��GOll�O|�1@l _�"�"XO��zHHTgϵ���k��K�c!{����8W!<aL���q�d���ҁ�چ�d���@����P��L:dQ�ˎ�&rt���t>U��k��ք�e7��:��Ë�^3�bM�;'B-��"C�a����cljhKt�>�D5'.M��o�J�8����Gs����� �K�%�.���.H^��#�Zim�u �?�y=m[}�o@����T�/�S>�����k�jo
���D�Q���}�)���P��X97����:A��[�c�-
�)K0����΋It�����E�C=��T���rsoU��b8ZD}!δ��y.�������c+q%T�h�;��{V����D��\�d�wcdy�]�?԰���1��*ϓv�]�>!������G�4=΃����Dj�MKFt %�-� svX��i��|3����T5I�P��c��(�{������6�U���x&Z�b��κ����Jppm��蛫C��HO.�T$w� %�5+���� �Y�h�'8�����$�⧠�O֝GO�SK��Y��ե	��B�o�p���U*�?۱B��,���6jX~���	["�%b�(4�1���J�ve�S��F�g�G�y�m��Q�:aI=��Z����7��#��� �ox��z%�������n�0F���Ѧ sڎ�N��c_a
�����c�N�])p��5���R�O˺"C׉eg���f4���(���lu�h	Zop��A`��F���a�>;�G#�����Ot�*Y��
���^.~,�D���w���ᚾ��u��>wgv	���/Z��69j0geaj>ƻ�gb�l`�Z��zg:hW��;^�uE�ʵ�f��v��X�K��T_5��Jh��]&܋
jEZm뛮�����vn��?����4^���E�WV��LIb���URQ)9�<�d�e�'�؎Fb*JY�91,H�o���#����k����.�^ȷ�X��'��8�A�	��m&�Ӟ�����6�� ��\�m�,�@
r����S��1�4�Ä�;��l1œ��*"d~�Y�9+V2�� ��G@���h��q������{_��#	�_��`4��:�)�>������
��dǏs��ҝ�DE�ňt}{�I�ܟ,��� t��	���)��蘇�4%n=����$�ߪ�C�:�넂z�ډi�N(�.�.���7�)�è��L��<n�1X��&�����Y?�_��pV��-������@�уai��f�ٙuc��J�DHJ:�^㲫7�6�IE/+�)/~ϙ>�T���e�Xu��;X��@���@���em�c������
�3��Bj�O�F(�w5�8����Y`O���|�I�t̕�����|����`F�mw�Wƒ+2N���Bl�]uL���n�ׯ;Z���SBe7�T6����H��B��q�'-#��˷�`<�찉�=��9�C}?$�k���}�~�M�,0����O6O����j���DH��F�u�?"�Ki���2��7MF�e�kj�V�9��=��֏����
��0��� 3{�E���g�m���;f�m���ā8��q3�&�٪���� �~�ﾘ���I˦�>�7���K\��'�-�Gi|�Ò"�ug*�rF	_,�NJ�(�TSQ�n�	��N�)Z=B�)Ȳ�w\�ө���]T�N���������(�[�j��J��H��Z�.��ہC�G���2bV�0@����FW�
#�P��}�/��tB���5-�7ri,?! 9-�A7FC�{?I��6/]�8,�K�I���Ԣ�y��q��(Ѡ��2v���	`�D4���q����Vm���
�+��=k�Y��gDm��
�ص�������Ǣ1.�� `Gd�n�;^�%���&䓋�|"�T�_��>*V�N6�X"�P���U��U�|��J�5�F�W{��ϤV�±��A�Ph�)z�����r��>���<V�9��&e���{]l6�1w�S�53���C|±H.i�f�S�48��t�x߸�������7�K��̨�|�`	RXc�S��C������[�I3�*���zƅ��T�8{*!�.Q���'��S_ �F��ג����*���� ��Q:��@�A��|
���X<�8��uo�MwF\-и?�>>�s墺*���O�7�0�b�3�B��`����(&�yp䯁��� pJaX<�lA�!.�<̌����UV��#2��pQ�ƎPQ�{Rw���.�A����%�"��e�%[��bf��5�lFҠ��kCWɺ+�)k~°ԫ��y��WK����r ^I���x��/xDO:f�e��9"�-�{� �x�H��|(<.�q6�GHy_��8��1��ɃWܸQ��8g�0��#?���a���e�#t��<��c��[B�p���p��� �%���W����YS�h��x���P*T!��>�~��q��{]�u ����4YtA�Z��Aׁe�	�8�dFi��� ��nT�j�����C��v�G�y��7����&?�C�3v?�7�#�+���L@���Ba�k	u�[�YV}�2Y���x��&�;ԡ!�ox���,p\�r�N�#{4��&�<e�Fo����5>��!�Q�0(��S֘=/�ոbP�����'�&�@v���'tB]�/m���&����@�8nZ��Y�ް�܌��%m3]S���޾ׂ���7�Pԥ,��%�\���5��=?!�Yy�U84+RÒ��p����B>G��(�HsuNH\,�I��Os����LBF���8ڢү�5�� l�)`�R\n/�X�Xy���'�1IF�C�u�B{X:P�TK�䙺� O
`Z��.�T@�x4(��o����ۥpӂ(0�y�ȸZ�'�뙥#�M����'��jԃ�nm2�w/��U��$�^˰I~%왯t��
:�*�'��`7����	��\%�oyn)���0�W�2����`��eZ��ܕ������R@@
�sg�O�G/�����ê��0��y:������X促��K��g,,ҥ0N�Oڒ��2E��X�B6{������"G+��4B��ӡW��Q�+,��k��^�
��Fg�Ѣ͜��3��Ƈ�w+K��{J/�A��MU~����b6�Nck��;��t����]$��m	;�u?��ڱ~N��
'���\P�ªK��Z?>�o=��x��愐P�,(�
����y�I�_�ְ�Ǆch�$�4ㄒ+�l��A���X�Gͧx4�o�EX� �r|�"|;*ϑ���j0�T}��Ƭ��,*tV�K�t{ȫ�����Q��e��b��8�&�@�Kְ�M��F�R܇���m]HN���P~��|��z�;�ԐC��n6D=��')�/`���#~S6M��dEk�OaL��+�4w�Q�%>�ae����E��]�^���K� �3��3*I���d��VxU���W�ʫ^%;�UnG)���u:�Hl������W�]R{�^~�XXP$���?��J6�e�iS�����{�|QA��]#���q`��q�5�i�$�}�������>^N�� @�UYe?&:m)=�;��2<��L�G�B!�&�C&j0�Rc�(�Y!	�~�i���:�On��\:]%�z�3�ٷ�_H�M�|����~̪��Za��8�d�+���d��5V�on��+��K8��l��:��GJ�{�	UִQ�e�m)e3~�x7�e��{% �������{�7|��~>b �_�	%&�%�sM=�\���}�x��Ҵ��C�*N��7ߚ*�H)�.&�2U��w��e_3ۚC�I07ק�&(eTD$5�ܯn�Vӿ�:㐓�����A��ss�ajU��'�q��8�/,v���4�9H�@8�:umw���u�?���:\�.��+�N3	!�+4��^�榟qr����L�]ʌ*�{�ePA�$oV��k$,�ʩ������2��<D�yj�k��ȳ8�����?���!&Mą�Q�����o��Cߌp.��`���ߨ�l�@%ۗ��$�Ko��2t���u�ܹ���vE�-�b�T�\�����$h�(!AG�j��0�B�A��O<��d�