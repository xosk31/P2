XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��%[C �@���ٷlO9e�;�?�G!���.� c��}-E���"��	��J�U-��[�}�HuҦ�Ig@��E_N9Q]��$�FM,0�Z��6�ӏ�*��V�c�x���d��`�޶�J+b���T�VDj:K�v����I�ʔ�S���q���)-� ��H�+S�E��P�	�J#�!A�d���Yv+%
L��׃s�1�H ��uk���z0���#<�PU����E)�,!]����4��2<��6u�Tk�oEn|� fN ��x��Q�=��,�rs�4���5� �h�d���(���ҬZ� �LbC�l� R*��d���*2JBx�H>MV��>�mO�-^�]� �y���^Ye��Y�K)����J�7�y���n�5��_O��������S$�o@�88�1־(��K�'?�9�}դȅd�t]�r$̠�~����
]`�9��If�4A5��� ز ��s�*���fϊ8d�eye�{Vd�pH�g��+!��7�aV�gm�C�����!���+�"vpæ>�٘HC�}�����l�M�,�I���t�*�\��6�z�ʀ`¿�1��-�#��o�h�ڡ�)��v|���j2*�6\۱{B�wa�����;%��L���������C46LCcd�%�q���	:��x��? �wTX==���%R?�Z��[F ,�����O�ݒ�-����-(a���ר�4ڒb�k=�p�D|��p]d~���J�C� �56��q�e'�2
�5
�z|Rf3��0�8XlxVHYEB    1e9e     910+���I��Ο#j8��������n,g�����ҁ�F3qSQ�z�_
��k,�ر9��G�39�v���F�~S�7�P�Bz|��g)*z��SDf�0W�NM�mNo�W�7��b��A�#��|7�W/�����2��4}����Y/fdO�vs���ApLޗ�O��ǉ�g&[m[4|f(��#B�9��A��1�����^�^:S�m������V���c�ܨr<K}�,��&�%�JcN���lR��*�kYb0C%�-2G�Gn*~{=~ ��������4��R'<��X'�d�>�x�볨��O�V�khу��eg�B;�A����R|@҈��|]X�����"be��B;�,6��b*�<b}�% A�߳�ֈ�S)���Л�^�R4���Ӡ�_:07�YLh��4w7���a�=����T�6m�����ns��<S�{����Y�Dty�Q� �
Og��NSI�>�`�֩��.�T@ш%ٷ���9!d�T�D�|���c��AS~2����{#��BC���"�yF�6BL�pt��r���b�33$^�1�1kǫ@�l�%���Q�8�*Lwj�,׌C��r$"�$J���)���k��?l�h���Q%= ��|�] �%t�~{D"��eg�6l,WYUx�>B>?8��kb��i� 9�f}�$+��h�.�3t��x��c�:���� ��z�s%�r�~������6"\�=�XB�ھꁟ<�k��:4�=���<��}=�p��R��5�����P�*�Φ�Z<��Tg�{,�9��Y�2 �b�?m}��ﾶ#��0xI����W_�g�;O���;�?̈́�����ID֦��:w5�;@8C�nN�H��k�z�%�NGgG���m�W�x��$�R����������,%sIsJ�ڸ������kBܢ	�N��h����U����1<6"�=��a�4�}ކj"�7�r�z׷� ���g?u����,�w#/,�mc���r�O��g7��W�u��dc�{��Sbi�9���g�a�"��Ə6��	/.^�]_��	�cn���WiO+�|����+���%r$�;�{�MՊ�$���vK/�{����YM��ఖ�C��"��r-��"��#���qo��>�ߑo4^�Va����'��梐si/71��~�5�K*sr��1�ic$�u<��Jm��!�6d���������o1��M���	�,[56Q��R��ܑ���Q7�,���'�-1��4�z��������C��xK	C�-����;���іi�cv7p� >v� �ƻV��� �ح�n�c6�3�m�ȝ����e������߿
�m�@@Y�*��`#�+
�蜀@�ð�{�I�C��\,�J�*��@_T9�^<�(�ϕ�D����[y�<qd����cc�~'i�1#�����9mz���؄��FD�&��iO��qm��_��|�D�l��5Y���:��Z��=&�Lp��]�C�XY9�7$��>�r
LQ?�F����!��ژ�9JhW@�⻣�iX�� ��0�m�mO��ImW�� ��m(�r瓷W�7���lo�Px��n�����k�2�L�n�\:���w~�i"a��X���(A�U�ߢq�IHк���c�kΜ���QkW�q�t	\��sJ�_Hv0�k5�
�dt�3A��|m���CZ�h=6��F<[a��Г܃z{j��j(p��Q�]�1B(>�E��4D�dp���BJŦy�2/�e~����_�uW=9�\=o�ڬ�.����0���ɬ�ē��=Dn��s��N��'�S�طb�5���D�������-Ίv�p�_K���Ć�O O�_byM��`2���������� �X���[��q����ċ2ncL���k*G#h��g2�>�7��q����X%��`YM����s8��v#��N�!��`3�n,=�?-�[���:E�eR�{�I�)�LZp=tB���u��DN1�Q:��h*�{٬��4��!� B����[�	���=����߳I0'��h�u.B�h*��,�8�Sڔm*4ʹ�&�Fؐr@�8�wf'"2��DPh�����sn�v�\�+�J��p`�_Q�+z_#��9�&�3�8j`˅W�B�Pݼ�u%H����۱��6��I�v��7s��;Gp�r�f8Y/+k���)��V��j�j��� �+���~��ޮ�5�S[3VT�!�݉|� �[B� �M�s~2���ܲ�xγ�N	�