XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��P�#�\'ap�z����e����4���,�J��qYE�v?�~�v}=��7)������Չl�푪+�2m���TjE��k4bk�)��N+ϓ-�s�1MY��b/�x���X��έ׍L=�e��{��V-��W�1��K��Ed�!�jٳ�,S�V;F<��ֹ����/sn�$+���`�[s��k�R����?U4�)����]�2_^��<�Jd����3<�����]�]0	�����I�L�����c�>�p�� �\�l'� p�������|��+3�J��@�:n�/c�?(��� ��������-0��b�M8Zˏ#���\��/8g�^�I�dU�����WBɝ�}]�KQ�<������D �M�w���㨬���UIkN��?����"���4�5��_;migw����2f�����NK�[@�w���k�C��By��a�gb��G4X��kLg�4�AӅ6��o>U��n8_�7xaSP݈n>e� �t�$ܢ���c��?�~z�-�k�/����e�A�B?�PV���f����"��ŠpQ�C�ӂ�K4g�95�_��N����<��Mnm��?�Wq��#�j�:�qb��<q��R�(�e8 �N�?6���d��*jL[�X �\9(�S�54����[3�L���ҡ�#��v#��ԍ�7u��j��@�9 6� 2�,�+�ɾH�.]����ʋu�O~��$�+����Ԟn���
������!}XlxVHYEB    fa00    2470�����Nyݜ��
�E�w�D�l9Kg��~��bC%�q�k���b���=��g��0eeJ� �`j+� %�I�S��&�
�b��-���{zIϗyК�0��^|��/�2�����`��D��b��;`[+X'J��J���~Դz)1�o�e@d�)(e�\���@�{@t���s#�4�>�t���k<���a�**��D�������-[�	<��t�t{M ��k k�!�J��v"��V^O) ���J�����ۊ"�F��P�N�4l� ��x`ہ�����\�쫉If񹀴. N�i=�S���6��� ��=�����VR��\�B�ߠ�N}&��R?]�.%8�$ʶR�����~�S�`s�#y��A���}8��{q'K���"��A��Z܎���5yrz���lߤ�
5�	wX�TH�����G
)�@�R��V��ɹ�(���6����k��u�d�}a1����3pC{�<��pE��kb�b�/�WRbkH��6,�����5s����ѿ�Ϻ߸0��!���dO�u��T����b�*�h%�R�^~����C�B�;� >-5N��#?�=�2� �>�����tQ5W3�m[z�kkg<�ߧ�2����q��:�6��F����@�t� CG۠��B��_	��Q���3�l�DE�����U�m��B*|�f�V��3t~5���.`�����|�����lɰ�o��`��V���{����&��#=ɰ��P{B���/_��VQ��v�=BO�_��o�Z\S5�n�w.:�ѽ��f��i��~�_��7�;���W�Z{�¹4�H�� l��:?�h�n"�ݡSs���V.��9n��+���H]�[HϜi����R�^mT�h�P%4}�����ڧ|4}��������n����qç~�gLT�f\����KfE-���!��?:�0����������g xA
����6��"|���3eP�S��c`j��q`��'���Q|?*�kY�H[���?���MȌ�����X(�?��R���d�,xz�1DᗸA���(�Vg`񣂞�Q�X� F"�T�h�+8�&�i�p\��2Kٻ�vds@��I=��Ǧ���3y&+=V��	9�b��xn5�p�����\���0����x�(���gi�	�=:` �-��
�Y��Pg�����wnN���9��*OFa���iE���1����
����́V$|\t���gQ�T1����]�%�ϵ���PR�6���T�Gk�?	<8�z�r�M���f��>\�O��<���d���!n#j�%�� �����R���8�΁��)�C2��������R�"95�Ij���]�٢:�ǁ�aة4O;�t]�wt%��� �C�w����ӂ��Wn�`�2��7�+V%B�:����fogX���(f��|�iGR�Jw$��s������Q�r�f�n��N�g2h��l�j'��	��|�b'�{~E V!�RC�Gv�E=5�/�H�69�9�Ӹ�+�y
ͫ����2�c��b����5A8��S=��{���m{����0PV��Ȕ�
���j`�1��	��5�{��a?'�5�����d&	Bei�I$�]��<�:S�o���r�j���3*&�Xt�A��A&�|y>����ig?@7�H]���>�;�X���Ȯ���ѥ�e|:J�_��s���eQ�OX����y���s�M�BT��oT��a"��6l4�қ�GK�?�?b��Zr��BeVK���8$Ɲ�v\�;����ŏ�#Y�u�c�c��������f<	�FVh�T�vZ3���[�Qv�Ĥ���yI���5����{�G��J�2�9��w��<q��w��c���:;�D�y����|���]�ȵrm&t$������Z	JJj��?U�Bo�0qV�9O�b��]��41isb�_��4��o��t^R`g��u(��<~�&��5Os��h!�wl��f����c5��b��;�ō�zy�d�iA9gtL ��6m?������'������B�E�>�7�!�ԗ�e��2�d���e��n�S��z�'���߃��voP@�Y==?Q��Df��t��2��qkO�(�w�qNaWv__{M��ǗM��O����w0���{x�3���������uX��0���+��L��ӎ�*�4����}� cQ��{L�f���rP�_u���z;�\o	M�[�]�PÀɃ�H�����XTΗU�Td)��uX*�\m�|@��@Ǣ(U�� w�#�i��\�YdD��ּR<5���]ju�#q^A�6�8��C�E�#�����V?�u�;�R� ~�p���L�ĳ���uF؄=0C��1��Ű�"�	N���,Pd�DL�� ��~�1�r�d�6����Q�	?y����yE�/K�q����L�*�tV�3��Y�yE�E���i�ë�DYaB ��b��78I��|r>���l���e�)��@�rI����Q>�ы��8o,�.Gr&��4�fw�'��d���&#��IQ�z���h�Cqk��%(��H܁���4�Y��);��^��#�ߨF���* )��G[�)h�Gv��s���у����(y��j-��T���mDL���JCk�"�(?1���B_�MŪ�B�h�6�l)3gw3��{{y�� ^2���Hp ��z����������_��q�z2�o��p��b���K��BIX�J�2�3�,��6���l�0%�����9"�1+�j���:� �P0T�AT�\�HVhg%���N��:����0v��b�ei�z�~��,�R�ܮ5�g��w ���Q�C��/�mvƈ�.,�P�E�؇K�47�lV�bI'�[J�!3Ut���"�P�|�Þ�ͨ��s{ic~����D��%@뱈:|�0� �h������N o7"�����~7C����]��X�I�^v�!��>�xC��R��ʆ�?{Z��m��^�f��!(u����������O�μ4��T�C-�-�)���܄�C�< ��-�jK�4l�l0OFf��Sv�~�+����u�A���WL�S�b�o�x0^ I����W;Ī����L�*RI�L��C���fP����� �� +O��)��-|�Tp;*�ͦ{�����4��y��%�;Á�&C���n�>a�cԍ����B@���|�v2-� ���z��\^^��!�m����o;xh����eIeUY�m ��4�h1���1�uk��	VW�%�O���nv�x��Zѥ��o���6na�Ȉ4���NY�������q`ŉ�5� 7���� �}ڽ���<WE����j�J���~���6Ҥ�x��D�'{+Y$-�����2��^2�ў֏�߹�B�}�ɗMc�z��\�4rq���]\Eg�F�,�EGm9����<\���A9M�$
�#�y�����T��Q����0z�}�L�P�n�Y�	��� ��A�y\�J���2`��fG_�^�T��3L�>%ה�ޣ�Uy��L�w���
i+'Z 9�/�}�d�����L��E��0�g�e���"i6")�t��2B�R��ٟ�0��M$*\�_�=��L��Q�Α)X���e�54a�uU���(k��Ő�%K4mD>�����7E�;��&m��(�,�D��~��4��F)�8s�������)�e�1��U+;���
/Ύd$6��ht�P3'%������j>�?�2I}�R�׈ٹx�9���J�I����@��W�":�a��e&uQU�.G���V���H(gKq��e�w/7�3I���<���-)�(����%O�J^<R��1�Ƴ�~�ns�w�G�ۈ���-��/�d�:k~-����zB������Wid�)>H��Yx���s�ڝ�36̙BQ<x���ڀ�����Ə�ϮpQu��'3.G���ep�t���%����!��s�����P\ÛI%3U=�>��ٝMQ#��F�cgJX68`���G�v�	L�Tq�]���3����j䑷�� Ip���s����So��/ၡn[ a�Qo����J5>�|�����? �@���U9���(�2��.�9@��p�M�0�M��0���N����>Ւ�h�M���j�F��6Bc24ߕ	�gp�tI	��V�����𡒵�����K�Q<��)��W�Xw|�]z�^�H�ߒ Y��
0���S˪����Je��4@.�uT�T�0X�[�WۍQ�{ťL�nY���o�D�l�Y~��8����ܘ2�de����FV��Z�oއ.n��=�-�Q�â�+)��O��.�MwftQ�Z&8���.(?KJ�w�W�%��3G�a+�^Z����f�._��hK��+�e=ɱj�����#��N܈�i�<{u*��$��<Ht-���ƴi��]K�K��������Y�[�1$�#��!ͦʠ�G��@h\�+7��|2��h#�NHs3P��D��vع��7�ȑ���ˀ>�@l��GBE)>�;��勘t�p�Q;���vs>�0��f)�;e��E��t��4{FFP����3�KE�^e�o~��UW�B����H��ʐ�tU>��ړk�k������Ŗ;�7&���\��G��!�;͵���+�K(!$p5�;5R(�W���+�='G3����CA�W����[�o�^80�W75��.Oq��N)�Tok�G:j]�]+��i"��7�!��{��Q)��г靴�PU���sF���=�3����71
����p*�je�M�"U7KD�)"�d_AOHk�vn�	�BQ� =6��Dʖsj2F�*ɻ�o|5�;I�J{�ǥp���<eݎ%���*{�?��'��G�_y&5ozUj��Cv���o�fo�#�po�6����8�Kb 1P,ɞ��%7�6�*��'�(�����o���05�ʍ�b�r:�񞃋=8ק���TȄ4�Ն����^�}����5EHa�rII-{l2>c�&{���߀GUlo������q�}.�wu�pylO�-��g'��=�����@(�G���4�/Ȅo�h��"�f�6�R���Ii�ޕ7��ԅ9o���$�	:��5����軉CS�}�.���<�:�h�j�SjJr�ج>ػj�W	}7J.����-�5F�����4u��䥱$h�-l�T���s;֨�Hp2M	�[�~�0��~�ѥ���J,���7IZ}�R���D��zCȝw�Jш�ū�RID��k��73"�X��.'Dti@6�����|.G�ܳ¸��>3l�P�:@[���\ժ��,L�l���s��Z���<!��-Tk��Ȫ�嶟)H�����E*��a*
K���s*g���Z�_v�a�����]']�_���닸��dz�����
A.��C��N���?�d�Mɞ�D2"J��dZ�CJ�rG#D��`��覫oK�+�w�^���㏻�{Έ�A"�+6S=T�o?m�nC�w%D���?{Y�����e���;�4�6�Z�����ZƎ$¡�o�]\Y2o���;�������>@��4<��%���o��c�BR����e���T ��q����OQwg^I/���J�v�Jj��DL%���b�B�L8�Y�S���[��_�����,��+hF���4��؝[r|�Cl"[��RF0뻌�z�s���t��O���B�8�«��'p�	��1����(R��{�K%�N(�S��Y���?k��.����ٔ���!թ)T���*��}^��[LFc[��W��9��ڋD�L������ ��!�c�D�qj��J��v������<=��	�](-��'�}a�f����M,P@S<V��pH[`1��tCB���P�@��\��ʦ��V^�Im���{����)�����X�,y_��f:/i�,b�Qi
��ۢ�Q�e�%�q�8��ᝑ1�c��~6Q���]2�^�%����L���6�" .����^�F)�p�+,����,�ߎ�:.ůZ��SK�t�_�(��@��a��T�z;��S��?��=���
�`	Z�â�l*3��+�/��O.�~�E˛�bk��8��C(4�z��V�ʢ,�5v�=������y����11*ϻ3gدv&uf-�����$��/�3F_!v�o��lpF��L]j\o	jUc���׽�,��q�iبR��	%�5�n
2z��&��<���p6�z��5��C�<P`Q�C79�O�m�Q��,�����Rٕ,%�����jvYd�r{b��>Ge��Ν�Lj4ο ;FH��.���ZP���35�3�,�4 �G��
���Zv*9���872Qt�s�\�fW���0q���x1��`b����G���$*xHj�,\�E����X�9��1F<��a�{FX�Ŀ��V��}7-�ͼ�p,iPVKxܠq	da���C}�F5�Z����[>֔f5����q�ukQ��e1��j._���L(U�:�fm��l>I����u����7?]A��3�DKr����"�v� ��)���Z_B�"{���c{��[�i!�D�b�OU�qo��K��W_��)��jӽ`W���h�P
F~�r�Lt4cw�~�"v��"uڸ����ʯ�W���`�����މm�'�a���m �/#��<�úsT�Yc�_��\��Q��bT8�_n	6���e'�G	�q@��K���@�ʋTjyw�Qb_�U�����7�c��@	lW@����T����5�ٲ����F�2۫��������VH1��"�K]����-�"���{����x�L�;�h��遽{Ȃ�ΛA���d��c�3���a��˶VC[*!�)މ��e�cv��w��(!c\
��2�~�Ht[�и/k)Q�����t�
�����2�&%<q�U&�5۴�Mv�!:l9j�>�ڈ=��~\����,I`Ӯ��D�he_��`յ�X��/�rF�8��"W������T��e�L�3��tq��:7E� Ū0��A���fi�N�T������u��D\��o��a��>,�pp�N�i'7,���4���v����1֠��V(jwNݕ�*�/��|���Mbj9���T��ZQ���C��Y:~\��ft�h���_oCW�d��)L �?se�S�sfN��vtz\���}V6�ҿ��;��b)���3��Ț�����B���6����
2ka��J̲��B�
�3���-����c=� w����ާc2�%fzrJ����r�N�H(;0��*�ט������gZ���ޱ{��Zɸ~)��m�q6������'������Yx�� \L�Gy�Az�.��"�!��\+�b7��oV�Ã�7���a�d޷����$�l�7/It�Q5(h�3XP%�I���~�#��h�u�^�p�M�=�����.Z-
�Rbﭡ�^T�����K����BQ��A�QÖf?Jܢ���Kw�ِ:�}�,�һ��ץ���u�`Ҍ�m=x�s�\��!9M��N����0��q ��%C�x7K����q�e@YT:�.[�OI%�0d�uN�H�k>�)�7yA��\g5�T��6]�۳���$�L<|4tX�+*��㰰S�OK�I/�¥HJ��4=�d����\H[w��V�+L�l�r�oJ��⌒܅�$�� ]Q<Qi��](c�^s� �(��	�����`=إ�]E.�P��c��$C�b��C���ik-U�dDhDb�Q�����[x��/e���N��M��w����MB�G��A��������'k{�)����V�}>�I|��6��u�R� �@�M<�e�zw[4�7>}����d�S��m��#��_��r]��P�����pgC��a��x�I�Z���6R��;N�M�K�Z�
#�*IO,�
�H�5���og�+������cNF�f'A� .5�bQҮ�D�Y�\��q��_��������)˼^�(�Y�M�8wQ�'�ه	���G贾�z�\y��hw+�v�ɖM�.�,�����H�r��=ߐ�[tm��H0��M�&�$���8�	�d
l���5;l�p.}���Ţj�P_�!T^O���2^��}Z��aѩ/秗��:������TRi����$��5�Hָw�B%=� A�\�~�\��AVx��atL�����	��h�[�	?MF'P���Q�t�Ze����P5��p�y�dCL^C���f�s�7;;K��!	��P�pL�m��;Ï(B~��$�g�a��<o���Jhڹ�7@wc��#i�!�V��ʄy�T+����}Š��F��%��.�Kn�[����;��%Ä��myf5���5�'/F:�����:�n�\�8��l���l���Y%�sc�������F�&yM�n��ǚ�i֊���X���&��0&��	�+Nc���}W~Ɋ��gש)�	�j6���R#:����1	�*
��p)Ǵ)T�kp�w����Iv�P����vk���y 詗*R1+�9z�=�c��ĕ�,2bP���S�q@Lcf����AyM)ƈ8N(��H���[����,H�X*-|I�xx��,��j)Ń+�t���k_�����i�!tQ�� S�4���xuVe���4��:�+���[������Es<8e2M��#�����.ጁ�%��v��ʗcܯ�+��n�D����� ����^Bu.�N�g�Z��:��C!N��K�Js��*1r��t��zBvnr��AGB�D^uf�� �*S(y�9��Z�6I/pJ`Mdލ��G����ȿb;Ԋ-*7������Ӂ�_ga�Z'g�����1'K��V�Vy�XW���B���-�j6��#�oR�Ggw$`&��<.v�iLi	�u����9�9(�Xzu����x�]�ʾ^���	J8�����
ݖ^�_(2d��������2���X�K��8!b�����*�޳�x"� AK�Y����8*߱�k�pf�T�=�#��5�R�GC��B�B�t�=�ԍ �`Me�#�^vnI�����y���s����ʩ���'��o��_�D�;Ӻי]�� n����
P�[i���#XlxVHYEB    fa00    1b30 �x��1BJ��t�����#p��Z.l-�=�40*Wt%��8�iP{0{لQ��,n4��_Rkh��ON���-���%��U�L�Ƞ2��,� �� ;��S������rk��0AR9��AU����הf�-����,?�p�7��j@a�%9 F���ܪ�t�U?uoo���P0xy�q0W�F֕�T�a��7z܍�sS&��XrA��
��q�6Z���0�>ɨa��d(�69G�\A�X6�=4~tm�:�qZ���]��<�$d ���B�1�{�`�SS��敊S��D�B��b����#�Uz�yOCfvejc�ڊل�1'�+�ς����t�Y!.�5{�q��T��T�7����-��lf�WYi�Dy�"���_[��^��c��(Y�'(�.�'be}�dAp� yӂ@�~��VW��\����ޮ�~�{^��� kJ��H!�{=$֚�P@`�et���+=uX�/�"`8C�^���0v����m��	�x.>��DN��� ��GX�R%k�L�J.i�B�y-�{��5j¦՘�I����-n�~ψ�[�nŧdW��d-.h)�)���N�I�t	�
t��&�J���j}���ϕ�2�m�k"E���<��ފ�H21Ro`���A�l_
-�(]�0�ةQ��)���m�j(���jm}�E�4B�jR����BRq-J�i+��EJh\'x<0�b@�t_O.6#,��&�ՓB�%��+ᘱ# �Id��?m���b&�����W�p/�VԞ;��9;U�)/@7�}�v*D$��Zr�}�!���k��&P�[���\��=�A���y�I���փы��b��2��!u����Ե6�N�䠿n�AO����b
�bMi�\�0'�ￇ�/�d���g�蔄;|�k�v�V��8�C��࿲%��8X<14J��'Y.�WU@��OW���Zw��a ���U�.����c^���#��S��ekm}ou��]�'�+�):Yj��I�2V�(����@Ma�E�c�;u�/T�
���M�o_�fO&�w�~]����_��ω�܏p�߬ jl���Z���э6������uָ��5%ĎҐg��|�q��������{^O�hc�;л��.&����K�>���qO �], C����@�;)�d��c�:�AoU��V���J��W��P)1�*��N߾��	B���mE�&��`j��1g�u����J7�2 W�T�^F}��.f�Bv�:�A�X��Qy�E[x�y�JR@�+�-k��ad�O,W�'��Sm��qK��/s>.�A��ǋt�t!w��F�J9�~%S��y�	NFxH�v�ʖ�.�Y	����I�	�j���1�G����I)��t���Q����b�t�L�v�8�WPr(�'q�n@���龬_��"j^�m��cJyG�U$�F"���=Z.��ѲԚuSi�Z�GA$ƚ�l�ݙ� >�nܸoM���W
�2��k{+��@*���@R����F��ۑM�8$87�<��P�HeW+��^�6&Ν(���X����8ҍ�Ԇ�l+�j�6�p����W��H��87���3�&\��v5W��0O1�����.|���N���ً�Ld؆���=��;ܲF�aJ�>~S�x�6x�����
�х{y6%)=��3mb�MN�X��h�9�QP��Y�`wJ��c��Lj����O�Lsi�`���Sԩ-ُ��H�ߓx	�Dˇ
Ɓ5�n\�Ti�S��Z���4� 	���k�[���K#A�w�\I�GN�#�'�ܰ���9ם3�"������xl�=�;-�[��2��(&EYT���f&2���-;]^֝S'�����=���r_��MoW�E~�����ںΊ�?H�}Ґ)�4��-�}ѫ��Z��ƵH�NxC���ib$g+��,��`m�S�M-Z�#�4��u�cM����W�^zfE�˺^�Цr���Ƀ@�HF�6��>4���[����{7hT`��Y��zr��N)��u�/�V Qyaj[�jwj��G�N$5�O6��,8�bّ��F�!�8˂-v
oD��Ȕ��.f�T$N�zVPA# 
_�d�)�Xx�i��w��� 9��zE�a�+��z`Ivq�k��*'
���C�۰�!J�0:ץ��C��0�A���"ێI��C{�<kMM��D�^�n�T���4Je�zc�f�T��p���Uў}�����`�14A��~�����H̍� ?��!}����r֕�0��##�/ǃ(���:�A;2_C�9.J8���k5�	������~ۙPI����=�tЪ�%���� �Zx�2�Nf����q�� �H6սV���+���D�/Zfc9oqf��j�"m^%��x��(���˅�1�����CPt?Ƅ�{_��	;F��zRm���(>2�^6 �uIL�iT�aɍQ7���?���](J6����m� ��5����[as��՟�:�a>&��pxi-:��:��C�ˬz{���V(更|��e]1�BpW]Z����Ȳmք���N2(j�q��c�J� P1<m���h�h�1x��~fU��=���e��E!i��4��ڄJ19�3j}�.bo
���N"�Q޹{�=ｱM��Μ"�P�;�&*;���h��� -Ѧ1�iQ��hx��>$U87&�D0+�R��,����&S�0K��q"7����l�U�����2�_������ȓ��v���������jD10�ˁ�Hق{X[�8լE嶾od��e>|�Z1�+�Ek�DW�$��'W����}�uH��ꛁ.�W�ĉ�����m�j��PΤcv�n���k���eŸO�7�޳�:���G�:��0���Qm�+E,K��|M[�rw;�2m�hC�� Q�@!d+V���X��KdjOgAx���Ӎ��[m�YFR{ �
�O�-Fh}΃�y�DDc<��l�:�j���?�=t0�Ч���ç\q�C�t8�:!�����:��]"H��$���	�;�>�{�֕g�/�4�E�A�8�#���ɱ��"�o��z��)��0R�wan٫��k��$�nF^���bD%�X��������6S8��c�v��g�n��oֿS�	��6*G���H$�Ix%�lE�H�p����H����fH%֠%�=0����;Jn� \h�ݳ��;69%a��M� q�6&	�� 0�����ˋ���]T�ɓ��IBt�F�;O�]f �\�p�s��[�<д<O!��-�vf
@�J���پc�����e؟�6t`�HE>�b�������_ {�!��R�>
;��Yr��6b'�q�Ⱥ����������-�Sop�a�L��D��j�@91�Ҹ�3w����S�pĠ��	>��$��&(5UD���bEr� kG�ۜ[k�P����snɃ�	����ϐ� k�/
�K��Ј-�Γ$�T�M+'�ǆ��~�dɢş���)Eqq�3��e;�
'N_k�)=v��M��w3��q�m�ʜ�6F�����Yw�� |5jK���;���Ī{w� V-�P�qb�r�\{����H���
����.�Y귯��� ���-^��vh�����\~�kŝ_�?�N�
�ό.
��f�O� y��f����0S{��!��9q��m,��[+� _���d�j�0��i�Z��~�{Ӄ0N�n�� s�?�Ht��Ĥd��}�k�#s�l�G�66:+�e:��ɹ���S7���-��!_�DT�՛c�l(A��H�59iR�m�������g}<�S�����b!����o����a�\��`�g�����	�m�V��0gD���0Qtv˯���"���� �3zaśEo�kUV ��^�6R�`W!�\
��/�M�70>i������Ϡ.�$�!��^�b 9*���@�m�,��zt���./om�&֭Y�j=�Tk�#���wK�g����PQ-2_� �u�Iԑ��n�0�����c�>��&I�s���ޙ)���b}���6�(fs��_��Rq`%�SW����o�<Ųn�)��7�u���2/�dsc8N��p*�q5�v6I�9�)6
b�eߊ�3�r�A8�sZ�|�(\sةC���wJÞQ٩�i��y��B�����G��5J^�hr��Uiz���W{
?�� �������\u�P5w,
�K�q���W�����4�jЄǭ<A�p�K��x���\iV�$�Y���Ċ/̔Qn�p��1H�C���C%�t7���Y|��V��ɞP��?��������_RY�a־���x��n� a���cs��8���Ta7gɇTٲhf���h��/
�p��1�E��ը��$��@�(���JnO	R�-2R�T��ݧ>:N;�x�5�-8��KF���t1�zlTۃ��YT�����E[�_xȳ��u��^Xʫ=�j�[�ښ2E0[Z�����S
l������\F<J�X-je�������Z�ï8y1�?G���U"Л�Sz�/�l�|�+�겾(��_�e�FT�T)���@J��mN�0��e���{��}ei^n��yu�p�pz�i��aN�%�^� ��s�K�@|x�.2�J��XBp{�5�OGR>�cݶK˻vy7�-�G鏽FO�/b��~`��sd%A�v�A�^����#}yid�Ivg�I=�|}��T1
��`�����Un:a�)�9��/�(^�ЋT	|�$W��,�z�����/��8�-CW���-DK�5�����[�+U�?_�$:���U���@+����k�����MtQ
�U����Y��+k��?ѤL[%��3L�8����pJw^����"�]�]K	��-Se׼9�n��N��s2Ut�ry m^��~�Gg�У�A,���_#'��t�>� ���}�d(j�n�d�Yy�7���e��X�S{�m{��4xr|x&i��f���2�mW7g5:��suiQ��Ed��^�r�l��ފ���k�3<�^sh�8Ú`oI���΍;	wy����.�Wb8���YV,�O��H��?�����41w��,ߕ�����	Y�b�ӦtHuX����t3V��ض7���2�2�"��2��^aZiK�s�\s��r�toԌ��NJ�����m���)Ա$��������@��h�T�g�0���d6S�q��N-�����TLE5�=՞�[Cy�����ku/?���OT��E��#2�L_̑G�}�m 3�I<�LH����Z��tW���x,�d	�� �"eF��h��m��g!�ܟ7�fA�gh�~���:�&���fQ��Oc=,�&��; /�aR�	�$,��[�Ԉ�����
&�4�6��5�{�*Ո?�N;�i�sr(j�>u�u�s�y	����1���/卵)N%�׭��`��� ��Z�͖#~�z�������~�5I�����������XJ����g�Qr���9-��d��ٮ��Uێ��ce��!����ުC��Y;r����@�F��)����g����g'��ucs|T�T�G��t�/�T+{�G��0� ҟ��+Z���ɐez�D.��t�<s�����df7��U��p��F,���/�+��="�j����:Q4}�|ݸ��&��I�i��⍲C���ޞ��{�v�df��Ǿ\W�y�r'� �6D�+�#�*���Ϧ�d�.����?AQ��X���������G#�g��
��b��F�"�T�yj���y��6���Z�X�~e���۟�h(2ŐKŔf	���ԤeX�>q����m1����k����wL!�ѐ�i�b�=�]5 ��`Gei���o�f����Ž{���MX�ۻ>	�[�V�����F���A"��\� li���\6Ȳ[O�3���w
�ZO���^m�����͑�5pLN+����b!��pv�ڹ�w!e�U^�<sPa'C �9�qA�ӑ~fc�+G�9�����G`i0?�1�
u�=�y�V��}��Щ����_ג�*��B�㴇��[2ԧ�+L�S�@��V�D��|���pRj�~``�Ἂ�,�e֤)+洜���u�B�$	t�)v}ADs�+>���s�����0��u'�>� �+��D^S�U\^����(��������5w��%9k�K_Wa�$���s�L��+3=���񙫹�i4�H�we"|1;��Q�tB{�Н*H�$��G��4������ul4j]`�蝙�>���%��1@���d[q�Z5w�:})վugx[��a!^n{)����t,eS}�dL�G	Y�8���Ѫ!��	��.�-��д�SԁR\�;V�_�:��m�Щ�����G���Sq�y���]d$�7#��S߰���l�X\'���|�
�:YwX����X.�զ@��Ewz;���\_$`�`�pz|�+4ڨa�@���3
�Ȥs��HVT�c���G�J���� !��~�r��O>W��bX���+L�/��b�;㱜@W�C�;�1��-�1hSѦ�#Zf��~��,5N��5mC�W^�U����./����J�1��mZ���.��j�EA�f��#���l�.AoI
�)�&&g`sW�it���b�I�Z��^�W{����)���cv��Qizn i��Xr;b��?V�3p�ɷ��R�*$�_�q���3��V��ww����T&7ϒ��S~5��QPƺ�׳U��WT`��1�nO؄�}��j�4g�J{�a�p~�˨�4]�ͻ� �k���AD}S��� �eݟ17�5�:���Gav@�V}�u�]�3l:=;��eX��CXlxVHYEB    fa00    1950(ʑsX�n�����vsY�e6�5���\)�Yj��seB
VbQSa�K��r�V����U�1E��6�S�1�j.� ���H�pd�/5M[�������� C��sڹ���Ӟ.w�-�$	�k[���h#������y���Կ�s��G�R������kI�&OP��%ڑN��-���t��s�D6�z���X��0�#d/_�x��ē��(%r�S�����U��]N���q�N��op#O�R
�l�#Go��W���V;$��e�pU+�%\�	Sy�����N!�b����p�ۄyA�J�ol�>��/�u�6X|�_�~JH�N֬?��\��%u�r%�lb��g@�m����0s3����;VV��0��y�,uœ*�D�a�*'2f�q5%���Q%�0�L�L}������@��.���41t"
��\4NgI�lY�$���GٽU�d���~H��!�UWY�+B���h�d���n"ν�L;@�&��3p��c��� ��]�K��Y�Ⲯ#olŕ�8����r%c�Q�\"�ÃI9R2�����f�k7��).�0�Cm������v��#��絭iv�o�����A��#����Y��vhRO�X@e�U�$'�F|�R[���H�����/�qF�bpCo���7�kT�y��[�Z݅|b�	BkJ��cꖾW7=
q"�X����/%�B��=���z�6]���/bes��}�J�0�����N{�l0hI��0>���tET=Bɷ�:h��d��9�<S���9G���� ���Y&rp�gl��Tt�wx���X Ю�.c����c9þQh�D�la�Aqv
h�&E��� ��l�z˰��y�#q�-ԥ���b�$ڹ1� -:5�k"D�͖�żߎ��o�:1�2���d����*�몴��0�&�N��T�䇉sܩɰv4$���>�1� 賧����"� $�m�v�(�#��'ݚ��	���55y%�����0���X�_^���n^���L��&$̷(��Rէ�?HH��┻�j�#��ᎉ1b�Aڲk�`�6?�B'�x"M8�H$4��%��6c���۪b	OvAϕ�q��)ay�XG��	2-VπJ3V������y�sĦ�3��AjY
^ �\���1���膯|{Y��a6���4�<.��{���Z���2�x'�'9�� ���˟�v���P;7~� �� �Ky]��t��pY��Y�Ax�`DB0����a1��GVXR\�������w݄El+��eT\�L~3_(n���Dq�h��X� dZ����ë*�G�<J뽪����Q%�� ]:�j�ĩ�n�ݶ�r,���`�� ��b���n��6��}�8b���m�D��We��h�������E8�r}��$��>�jP	�nW��Ny��V���!����f@o�!�7�{7��x\���v���Z����rj���Z*�jKj�%��ҧ���0z	�����ؒ�5��h�.�{���c��'q�I�"v[��������ߨ��g� ޑBʄq��`*���3A�j:���>��@�.]��;��@��q���[��[]�I@Kψ�]�h9�L�e�{� 7㣮q�e3\�R ƃ!��*���B��9@`��G�������%G��s�r��ƧI�7��I��I�k�=0gw{���v�~�z�K�5+[N-�c�r���㔱J�Z�ǎ��EGzlw��F�86Ѿ����'l^�*W�M)��a3Q���tK�$ ����7������w)�!����AT��5ϊ|���$OΌ/���' )�@�7�=����E~���b?�������k�S��r���#+|�{�"|"�K�'��_É)�Y�D/CG�\DT�_0і�+�h+���A� 5(2�q3��z�޺#������I����uW?�e��1�~:ǎɷ=�r4�>�������q�A椖vE�fC�P�Lz�Ļ�Z�����[�.�,#�CX�+A`K� �
��1���P��,
�`匕�f������s �&^Aw�ˌ����^$�1ӝ���L3���6>r
;[.t���).�ϹF�����ϸj�}^LS��ײ �a�Y��E0B����D��5���ܺ�����})_!�7Qq�SF�8���dK��H�>�X�i���j���B.��B��nAY��m`���yy[��d���v{(�0F�	M6�Z#�J6n[nN�HЯ�?�K[�?a��EX��H�+h'�"V�Rx1�Q�Fbeд��j-�%G����h�9�#{��i�Ԕ���1��'Nf��}Ič�Y59L%����N�z�S���$�Uu�A���`ޫ��΋���kh~P�K���w�O��uW� ����ǞP?�.�ۄ#*"`7:+�B�����9���?�^����������c�e��= �:(�A�5gO>�H��N4s���@�{��׏W4��f7/āxvv�H�Rs�/����֘�災���Qn_����zc�|B����R�!e�1�u�T�WEk ��A��o��,>�Y^V�����b��z
>����ԽӾ�T���-����6/��{��1T
��)=BV���+�2�-XZ�6�'}�A̷KV=�Jd���'���
a�2Ai��E���`��V�k[�:9��]�H���FN�E#J�hJi�oѤ�,j%N����3�%�"��Mq�\��+Ɏ��\�D��(��f�E����z����g*9��"��y�Xf0%���͐[t��3$�]NA��I�47�@��B�L�pN<�n���:QHx�;�����(�r�쉵Aզ�,�s`mPDrX�D����+�S�bz<ru�x���Bȉ4׶W�;f�Jr�VY���Nb�)�\�>�^�x��/6�^���º����GH=��i��v�
D5�t-9��j '���3Db�*[�S�_a �H<x��.T��_��s�$�*�����S�DTuM�`)�Gξb�[�������	��j�Z�����ªrs���-V8D��&L�g?���2K ��d!�S宿��d^id�	�����O5��x.<�|����Ah�����*uZ¬ܫOR�B��cZ�m1W5���<�eQ��$�hAi+�g���
k�>AL�ݲ���,w��g�%�(x�ćb�iͤ�9D9�����T��ט�P����U#���[Y^'*��)m_�(f�z9˯D|oþ��Z;�;/�+�	hՀ�}f��jE�t�:�p�؄da�Viz������s�����n�)���3�2t�`2|w�3R��C0�j���h��O�|C 	}M��ƽ昇v�OP�D���B�ݖ��L�,0E��{�O\��c7mNy�E!v�j�Pli<� J��>���9��2�o
 ,��k�K%w�!��^�"H�:'�#S���@M���q:�t�-��M�"�Q>��Q	�b��55���ww�dLg$M�aN�������M��>sZ��.��!�Z��mB�ҖgP����mf��(z9?���t��ܬ^�E�D,�?�ذ�L���|0;�f/����g>�����os��$���Ӕ:2̷'/t��m�r�	NG�%�QY��=#���ي��x��Цq��0B��w[�%�=+ �/k��~32G�/+ilʗ�^�]ZK�ݟB�� ������w���	��]yJ�Khv*���������~�Wm�Ql��%�u�h�	�YV���L�)+J��P�&O#����+��9�������m�3�d?.~�ioD�@�B�1O�<H��2�P6�Y K�X��bȭ��`����?Z+Cҋ���WY�͘/2-z�h\�_v�L�O����)v��_0fa�6|�4�it	9K�xg���{l`�����z����B�~D�xH���L�,y�*^����F(B���T�^l�Ȅ��5Ά�-� Zw,��H�
�}u�����p��b�}]�O��B�5_eLdЀu��4�7���ji��q��7f�O^���B���a��y.��aW��u'���Fl5�ӊ�L��=uf)��U��2/w^�'g�\-�b3H�=[�_��k�E.�u�z4��d�%	ws3��!~*�����J8�Xq�<�2tO
���Y��pt�w�)���N��e�N�a4���<�s�~dS��%��qҩ��Y]�@U�۠c�g� �ң#)$�(,оX�#~�����
q��f��J.37l-b��R������D2v�'�?����7 g�f�:y$�χ2Y��Ldώ���A�L��S0���j�
B}��$t�]�M��i�12:�~L��&�D�e'#ɃP.r��(�!��PN�I(W?�&�Po%��d�&�*&�3A�/� ���_�@�c�R����f��#?`��Y��-��ˎ��7+w"#����υov�UP&�B?�a�Wѿ��Gh������tc3���e�.�Rv����£��PZ���-<E�w��cטnG�A?�PN��_�˱우h�?3F,�����.7p��v�H"��=X���-�2�4֍䪄��P��t>ԅ0�`�6(���2Q�������/`@��3��̰ҍ��9w�;�@dE[���)j��Y�.��BP]R)v��d��#x�z�@��D�C%���Zػ�qU� ��7��;c��;e<ﾔ��據��L����]o�A�aK�d:��_���Iv<��pY�Nc�K�ܶ��o#x^�Q���Er��5f�,��ɮ���� ���X���z��g"�W���H��b,����F�i�&��oI�C9\8�/�~�|%�e+i@ B�2��fMÌ"��2?5�G�p��+c���6.��Q�B][�����QZ��ee�����(O�i������P�U�	������u��&�����oDכ*'S;��`*�� ]p��C���&�n`�����}�*���Ѻ��u�U˺/9f!̋º�o"�?����V���ڴ��%�q��V|�0{)=��6�ΐ��(�S��}H��[�6�9�bP3�R���&z�R ����G��i�j�hW֯s$����[�����64�w+��jQg�s��ov�.n�
�C^�K����<IF� 2�׈�`8x̖��o�E�s���]�3
����2k]��2��hL�v�3�d��SX�d���d�KԬsR�!�v������˩*�'
G鐓7��7
��#����-zb�r%���l�w���:���fwF��E��I�ir�J�v����$7"��U��)���烾5��q�xsU�P��G�89��0׈��v ��X� �}П=6v-X��q��\s1��P(#?�ȍ��iO�ȗ�\��&�w{P;��$�<&Ay��� ����_-�� EQ���1^-�?b�M":�)@�<�0���������o�c��K�q�;̓��j�ib�ƍ>u�E�z������MeN �����B��R��������FX��V��#��u5������_j��{A�p��}V"�Ɯ��qpX����Z�q�Kz�k���R{bm+'��{%�����f�g�?��tzL�e����Hpq���sX2��^����i��tR�^���z��Bs�r��?g�p�j��u�,hgٴR��ҫ1}ot0�c{���M��gy�Ht�o����0s���c����JD$�U!&N�#���]{v�=�%�/�g���������Z?<d.��Ő'03Qr�iw�S��pb ��)z��Ȃ��j!��5g�����6�K|0$�@;��Y�c���Z�u�/���{VI�<A5��S�Q0���Ҽ|�j����Ff����I��2�:>ن�0ӽ��!~	Ex��KS��g��%�s��ߦ��Tc�3�辌*�z��)]]P�̕�c�د�6�50��0R@M��O&0�� �x�c�{�f��G��SYna�ıَ!�k٩�r����Ћ�-F�HN�>s!��9������1=��g>�� ���Ѕ�z;]��m�9��v#d�Y�i�����D�����[�a�گop�l3�n<�-������"�����]ō�{Xi�"�������ǗN��+X���u�1�[-Q�Y�L�#�����j;�/��md�[�_`�nq���z��fs�T�U��Y�r�6��"D�5����[>�������f�[�[\k̉���HJ;8x9s�?���=s��j��_�=���o	����$�gé�@�+:�S��B�H���VEP�x"i�t`졋�.e���}����̅K�QX�e+�@���5����%�!y�[,��XlxVHYEB    4f27     d40�U���ב���RT��`
�oS�ܢ�L���?�{�����C%<�	
���#��;�\���U��詑�V�=z��B�4��sP���5���z�t)&vp����O���̓��O͠zxcU~�}���#(>9�mn���.�sb��	�����:(��jaҗ��I�]lm�8ș5��ļ�+M�_g��S�M~�{�A�p�΀�w��X�}G�� ��}Kw��t�x���B�ru:�	9s���.+2�1�%�Q�9�D���4��+z�`�`�P�M#��K'�sdR>�@h��7���v\�����R��kJ@v��o|��_<�sP4�SF�14X��-QC��_@'�r�V�#�|��|��Z��s�p;��+���p뼉�%�uƄ�m��S-�Y�͵���HE'��8 m2��h�l��&A�ڂ�]�գٲG��6��#;��c�ڡ�s�n�3�R>��^]�{�{q�R+�H�^��?�Q�d>������B4�2}��N�0��T��	w��<��C��Kmg��EQ^SO> (�8�ǒGMs��e�q>��~�$�����98t�=P��PVR��s0�D�uKv��g�<J����w�U�3��j��Þ�y��%�yE����TG3�%�%qޗ�dy��; �e��p0,\dc�O �ñ�=���+B�K&vبw�*a�XOҗS�m�c����u7h �Ǭ���~_C�7��^�U]_��|�聱��m�>"-]�f'	���J���Y��Y�9��M���'��%�#�R�ˉ�&�������"�Cf���X�8oRr��j�7�����u)�S?�����z\��N�6�%�sP9���! ������\�_q�-
��F�r&{��Y�"Mj�D\�[LK�l��5=�?��,h��X{˾�43`/�m�%��T9Ï*^��g�n�2�o��I���)��m��ÔP���0��J	�_s�gV.�[�0��/���QiBBG��{$��,M!p��{W��*��9���3Cn�cMHH�诃s�k��~����:��<��W��`��Q{�����M�ȁ�6�@�3�r.��.�Q�K���1�*�ۚ6t�������!_�e�=f���|�I���r��h����/�mz� �=c`&ʹ�5�ktԶ(������W��x+."a���h�o����VUR��Bs1k��a�Os�},��80�T�����,X��vc���F��!��I�� �a�UI��H�M�OO�9�� ��#�L���fT�^P��K���~��j�q��ܱ��,��Q�-�|��ِӒ������)��PmCts��m�`|]��v,���7EY��?׍cN��6�b�n��)|ӏx[�{X�lV��"�+BָX��ǉ�L��2��M_rR�F��Щ���"ⒺW�˅��p�|wr�u)�F�����ɼ�n�|�)�Vw�+�����8�R臽�|��5Bш,�K����" ~w*�&�*�����].J�Lj��GwT����w]a����2\b�Q��i�q?�/p���4v�K���Y����c��$l�_8����?�'�s���pֺ��������plf=���gy�;�6�w����]�9^�����}�q�FZ�ؒ�c`&Rm3}�sQ�vR	���r�A��ϋ���.:C���<v%������?�Ƞ���\�lEoj;���D�6��h���_��i�n�u��9�ÍYrß0��#) ��n&#��T4����d�D��!�u��;��'�*N���(go�n߅�m{[X#}�7������B��¸�]�6f�nW�+��1D�.�f���i��<��<�xԻy�i� +���T����Q�ʱI{m�"� J_�gp�]�����s�c�ɬWp�J�#�33��.�6a�El�9*��E���Ԑ(!n9�ϲ"W��~7PY/���Qݵ������Y�dklDc���+�Cޣj��7�/������@����p{]������oL����ơ��u����
URdn�P]μ<7��Oz�${8��㺢;���f�4���;����'n�ǆK�b�溦$��:Q{O�WD�RI�Cs)+%�ާu����ӓ^ܷ�\��;�e�,�j��3�b�y�Jt\�PE�KP; A�(j�� ژJ�����}d{����X�=�Os�%�M�����< ��6.��ǺW�(X�<T�Z｠�p(�ʕ�_��r�-Q�KM���DQ݌�ئ��m���p��O!aU�!���o�T���IHѭ�sKz7��Sj/q���u'�]�e��(���
۩��Sk�P��j�[�k���엒��Oq�����|4���`q-�I\D�٧���M�H��#�*�$�\Q��F���ކP&5V_���n�~ʳ�ޛ�,���<�p!RXS�ӅKُ�\�2�_�-x��,��:��Ey�FIT�=��H���BNP��b_--M|�@�yF�o�xe�i[��Ϫ�������"̨�}��۵!��f���:��s#W��12���}X�U����3B¸XQ�L��Q3x�e�N
�R6l�27�v���W����tk	8����J�WK��<��8u2F;�Ͳ�����l��Ǐ�2��*��?x��H���₁'NQ
Ş{4'�p=g�y��f��J���Gi��q���c�EL:X�[p| ��n�F�"x����i�9I�{QlH�&V��F���#���đ)ai������m���˹ +���1�ƾ�|!4��Ì�����*/�Hs&�8rTč�0=�`�x��?(-�˗3;Mey;�L� }�s�K�U��sMW����'��U'�[Y����7���;��Ty4v����`Ӥmw���ju0D-�3�ª�p/�ܻ�����cAN��c}0�\R��8M��ݗ;��耛�i�5�/947;)�֜f�����|$Q��)�<���G�v^�n}.s 0����������T9P�j����S�?���C�"Փ���)s��r-�ޗ�x)�Ӿ�B����Dtx1'��lD}�7J"
�;1������]3V�@�����A 9+���/a%��^gJl�z��|q"�Ŭ�f�7GCZP�\�k�%�s�ܛnhS�7��G*�f����;�v���H.���?�n�d�R�����\�`G�c��=76"x�8S*�$��R�\G�Q2�}��%3��8�
�$)IȔ���������!o�Z�������GE�f���w��֖�(�4�#?r����<�GofKi���U+