XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����ٽVO�wn4s�!zp�,@T�i����V��w�R pe@�(=̤�rFib.���8�ȇ��8eC���n�R�2�ӋuD�<�Ҥx�ǼU7.j.}��FKQ!�j��Lv`�q*X$-V��<��C[7�fGlq6=�{�L�����O�]"�ƴ�͖&;�#GAN���Dh-Edt�u�U+�Lܞ��<����UV�iy���m:ץ��z�qv�X{6bpd���(+CB�����������>JS�7ɡ�V���ɟf&�̇D�~�f�kRr���X�chha���IK/�x�@�o~I�Pn���L�G�~�x7��Ͽ��9W�ɮ3���"���#7�R��aĳ/t�"W������ʗ��K��if�����"=x�T�F�	�Mȇ �%#]��fp��3V	����ū��('�ڔND�r����v.�*���=���t�e]|�[L���L���*xD�-qg���!�_W��n�P�SIw��42{{��].(�~����4um0�y��'�
�	a�v����'M�F �*L��u(�Q&@8�����T>��m��0{G����I�v\Ά�9��K�7ZR�)V>H���qw�ѕ2�D��<N�ӎn��>��>�@���7��zo�R��VHDK!��-x✧�&��ߙ�>ͦWAjݗ�H�|�Ly�c�`(����=�+��?�	)��*Zf��=�	�l���t��sqh�g1��x���(ZG��1|T���@�ܜ.ކ��[1�!?Ѯ�XlxVHYEB    1aef     9503�^�Pj3����P�7�A�M��k �D�][��\�r��
����C.�׼��%L�����S��,��V��1����V&^\�g�(I��<��~�S��t��uM��I]�D_��3��<@M��[\���:(������A0ntD����@l����ͱ�j!;ԯ�ʕ�:�_ے�k1�;��%t2��1w�"�&o<HkR��_��2�
(Ӽ[[]3h�h{W[9�ݎ�t�5M�q��Mnd7K�b/}-�#�K��1��3�Y۶�:�j�M������i� U練(߾�zO`��;n�pW��G�	��:�Wm���\hF6�����	��IB&M�<�̸m���3��6��,����U4�|������قc�m�������b�ҹ���d r!	�s>G� ��}�������a:��5ƒ<�G)}qXAA�V�_D�c"������q	Үʁk��pk���3�TyFlOɮF�A��������z� ��	5lCU��D�8/D5���i��.r�s�p��k}G(I���3�l�ũ��q�"�����+��0����b��0��iʵ���H�E��@=��y��m�e��s��4�����6�k�W`��b�2�&�DI�4�ef)E��)��ڍ
���%�+2�t�uP�cp��YZ@�θ V�����.g���]?�pՃ5YQ�Bm�@��V���O&�l��,  Ykk�[�&^�Y��i���%u�Fs,ZJ�ƽk!��R���k�:�����c����`ū�a����o�)�C6 �Զ��b+���[�o�^��,�j���Ƭ�Վ��_ϠODa?�0��h�q�Jb�����-"���ߖ�t.5o�}פ�O�Ń[�Gw���p���o��m�	`<�|�4����0�/�Ѕ�1�r��q�^�Rn&����ז�������l����S �B<�ud�k��@��_ٿjIU΃�� �������S�r=��4@�.5�P��8���9�H�`�<�N�-�t� ���
Ck��+�yރ��Ӈsٱ����F�a����[�)#��P���<W|�H8��1�w��/�'��&���b>�� �_��s�LNCb	l��vZ5�&�!��k<:S���ݽ�!���E)6������E��iͦ(x7��C=��G�/�

'4�c[0!(eL��-v���{Q,�Ǿ���C��R�XP�ēG���U	��ØZ�����9H3ۜu��Z.�''8��r'����d�-������Z�x�\�������[��x!W,�v%�x�ĶG����J�G��_���<�i�gcLcqBs;a���wo	��c�	��s�U�:�V��%���@��0;z�u|e��hB]~1\�w���!Vn��������5%��9T9~q�spȖ>�-I�d2ѫ�� j!�{�3���0�l�jr8���YN"y�qTkN�9�tzO��:�)�S�d���G�r��+oF݋�{�mp(��4���|r5��n����qV�ZI� Σ�m��U�Q��׬��d��%<_�I��'#T,DAy(�o�aM��wc #7!�!��̦����|����7s7
5��d��ST���S�Z9]��Cn����zH
��1J>�J߶A�(s��w���Ꞩ��r�A��S�Fu6<q�\&�0k2?�	�@�x=wż�@`gW�IB��uOM��K,�򤝤`�x
��i��-���������E,2��o��\p~����+G�+x�q��f�=���б�u0G^�";I�!3f����h�塎X�!xnh!,u�ޯ�G~g� ��\6lc)DV��N'a��zTn��������ۅ����x�]lX��
a8ʠ�-s
xb�qfj&���g�`�h��v����t#�[�s��Y��^�Љɏfc�pWV��=6.�\�Q����/9���a��e�́�>h��kQ= bnٜ0Y����'8��!����ٺ�`'�,�����8[�W��M'5#I�uM���[��z'���+��e�.�|��ZtT��m��	�����myo#ﵯ_
�?Iq3���BF���<����>�4,��w���3QN���:(K�i�^����rWW�1���J���@f#w��D�Y19k�!�K��#� c躰8�MV,mړ7���6�X��+�iA�%����|�zkA,��,ua;��0}��Wɛ!v�Dw�W���Qb��{S�z�87܅7��ܖ���I:ͼyꀀKQ���2`\u���Z��Ov1&ˬ]��#��kƏ�}��6�5>r��'�������@xJj��Q�v�񧚀Ҿ