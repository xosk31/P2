XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����h�!�P��2�X�5\��ʩu��ME���9�����}� y	g������2�f�
�yI�~�����)ߊ���������\�S��D�5�A"B-�yɰ�귍�I3��q^:w;>tǳ 4<3��۞�}P�8~J��x�Lߧ:�V��0��5��e~u��F��f��U\�*���GB�wA�=��\6�{c���K�n��1�nȃ��]h*oB {乘���[����h��2��~�q�A͖��۸;��@\!7$���QLժ�T�l����3j����;	H<�i�Cb���b���Q\�𶵏�xY��BL#>�[�|�$�R���B�� vW����>3mɘs�+�Tc}K�.Y���P'
��p�VS��
`���J ����uт
��7j5�רU%�3�5i��c�/�j��k�L<��B��K��|���
��Y�O�R�y�h�fb�Yu�����@t��������o2��:\�&����>��p�J��^@�B_����ow³�Tq0�~/�D�K�s���\O*%������҆��K����u�"چ8�6�����9%����6����		���чٟ��/�W���{k!��Z��w�����f����E"��K'�Y��a��6�%�]�`&c0~>��.>Yb0`GG2\��	����	�eQ\ ����ש���Лo�����П�j��u���<����]U����:w����
�	�`�H��i�r�7��r�<�bx�wbؒXlxVHYEB    1ce4     9e0#�gz���^*9D�o�z�)��< +�x�'��������4|;Yǈ���u}�l6�9����v�DS�G�p������V>f�9j�=}�u�1˳��7n�Bo����5V��G��.е*8�$����H�������L�5b6����u����r�ޓ�]S��S�@l�O��Ԝ�s�>��I�ȶ�/7G��/
{<]^���~�LUD������w�q!���R9Q@p�$�G:[V�o߆�����SFe�t4�&ش��i����!�t
���ܽ^�|�������$E����Ls�X!��D�'���f����`2S�\��܄�A�AJt�]�O��Y�Q�Xh���2r�O��~c ������/u�#�ocx��MF�褷�UN�,�M��S���.�+�>�+:Bo[�<�s�����&��������
���33'��%�?��ȩ}���R�8�)�P�����}�-�'3 �k/y׳ ϯ��쯵�_�H�/jC#�^v�2�cJ��-�qk@#�
C�(C������5Ě��F���,OƮZPl�c9\��f��\6�|�T�*��^Ϫ�,P�Gi߀_Ʋ蹪Mu�h�&���!3�����q� �(�z(�_���~Nu¥�)��~O�y���-'֔BA�P0!{���V��3���Ul�s���k���I@�P>㠳gQy�$�5���G|05E��S�P�j1�B[��\��kD�K�7��6%A�YK�ř�?�;�B\�^_��\~If�,AVr���5U�4}kC,.m�s��xo�͋ ��nh3Z�cX�-['F�W�l���x|�\rH#7�{Zg��b-s�R0���8R� �_��P+��v�e��3����&ϷO�i�C�u��q����+X��AM���G�-��g�݂w1���αj�lO)�w��>�bt��WC1����тUK��h�4��g�{,��"u��P�Ó�nVc��o�����kק(k��1���%�s��g�"�������|5+װ�pʳ����a~�氄�;���dx�h��������3|�ܯ�5�X��*�$����F?���� :r���_`x�ef"�C��=�^-Up�M�T���\4�Ί���[O`��!�uKCy�TB<l4l�r����n���q
�Z�$!r%�4�r�u�| ���xR4V6�jz��(6ȥ	���13N��fN#���~[3����zz�t*d
���k���25杏{Pk�w�c�O��&k3ǣFax*oj�o���u�iQ}���<�{~��v��'������=T�"8�f�b��W���o�g���=3B���ʒ�d������d�M���U���з���h��ܬPb�a�cM��B��ٽ&��P�I��2�������n�u��
۷f �#��f�t�xje�2�S�1��;FP�ZNᧆ�:���i��-�cWM6�%�S@8'�)4B����C��|��uK���@L��
�bӣ&{�n<5s�c���/}�#�*V�K�݂�$�������;F�/�3L�tF~X;_��痮���~�>[2G!���ȭ�yu1(3�)8��Zˁ�����^�����ͽ���9��k?/V�X�Ӽ������ƴ�����c�w�
�I5���+7�Ϯ��.�p4[�S�/`2p��#f��X�هA��42t�Lnk���&v쀩�JE��7n������I@�Ws�r��ށ)Bu?�{u��L��e'�-nK5R*�K�y.�җA� @�Q\uN�ej�t�����"�Ю� �掞��p���N����۔d��8�	�x3��������췭M%���P.��`�X*�V����z��~�n��~ȋ>Y"#	T���^���QR�@�n�L��Z�:�{��]u@�"nt�S�����W�qT8�j��1�I'C�T��O�i��ҲUk�mb��rZ�;��@jp>�!hI��~�4�b�ժxW��Wr��SoU�cVm�Jt�H�����]�*D�����q*��z�ɧrY��3߅��F2�e�Ɋ �L�� T(���p��o"s�)H�4}9^(���f����C:�O�=����Ե� ���� �^e%�.�h��ŕ�#u�|�xm!I�LB�d����^����ST�[�w��wg�O7��0��/vJ�����Z�ޚ�r��{�&ô��oX�0�t5@[��7=�Q��m:����|]Y�S�0��r�EB��$� �d��Ϛ������\��`�P��T�7��t"���B�ÿ0��vGJQ��i�9x�^�.��}��CF5��� �Ԓ0�~��G��6��ړ�Wi�j,u��ժr��uQ�w�c�{r<6V���Q_�����j��/a�'�_���MF�:��Þ�%�8���z�E�j�߄oC��%�@�䯱_x�n�H�+)����?�[�Ui�5�r�M��H͍+7��	