XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���+���M��N�G�`<c�y��C�E���q;�O�����f��Mw�V����o�{��By�l\G�$˟#�����w���[Л)^���{mk.K���ۊ�G�
���}����w�Z�O���"�����d��f�	R��?��p��A׼mI�j?�%"i�"]I5�x��{5J��"Q+�z�c������4���U������P���t�>�E�d�Pi����Gn����>�  ^-Cz�^�.���'�v�������=�H���.�"�c�^�z�G.��6F�
cĲ��P���̪�0�DL�Ъ�����ي9����[����dܒ���� U����H��)�0��0 �,�9�G��:l���K>�!����Ȏ^�������+)^J$�7-ͽF3Jc?���1^����k��OM�q�0�D�v�qlЕU3t��i�I ����qoؓژ�{h�)��ԫn�־���LT�}ٯ��m��=���*5|����3��w��ň��]~�o�'��b�3���C��˕�����6[�/a$���'W��K<��R�f�d�SQT.!}��><����0�|	�
[2�U�)�d2%����-�!뙍���R�C(��Ut��~'��̗܀9��B���p딳�^N���V��ih"���U!��n���7��l�s���`]�l���v��i #�D���ȶY��Ϗ�
�R���/�&	E]M�-��<��t�x�,��ɴ0�@ڼ��#�']H�XlxVHYEB    1da6     940kbo�^�k<D��MaM�QÜ�d���CMs�亠$�1��!-�H�i�AM���.d#
�x��w��*G��0�ٖH7�p���_�-J.�1	 ʈ�N�
���W*�Xܲ��7�^ZQ����@|�'۹2�p���-�;���E��r�1!sS(޳m&���~��i	][]hi\�Ti�>���P�wͤ[D��5�>�z\R���4�d���	�"L�P�+� ����MU��`��\6)
����T�RE~����X�a 	\��ų���IZ��z��*ժnH]7����q��M���rOq�!��V�}K0v�������cZ�K�L��w'��fmo��{�%��U䊹�~{�8D��r�d�Dt�&� ۗl�5�~�Ur�6���EEſ�b��,e-� ���y���H���:�_N������%���e���[^��)~���l&g>*5�?C^thr�����Ԩ`�';�.�脍c�N���\������S���@���(���f���v�,|"�t>��PTJ~���V�+;���Dzx�'���À ��#F����v�RP�	4KWS��Eߍҍ��&�/6��)��6jȱx�<���{+�3�^g��
_t���B�<k�[r��I�d��p+
»Ѻ���W4�ߎ��.!�&ՠ��B}iM},n��X0�O��h�t=5bya��)�Q�q���z���/n�b�\�F����<�hM^������&�tCB���"8.�p��+0������\���@�=bJ������!n������� ��7�^��]i�7��H�ǥQ5c��~��MN�u��yF��U"&�I�}�U.�N���5��	{a��yx��1ΨqIS�g�����
~����;;(�[ٻ�^�="��
X���0�Z�	 ��^)�
��6P ��3�r��`��O�eE�l��ۙ��z`�/a���(��f�������FLf��;ts�3ǚ�6G�����xd����	ɇ>��eLVG��y�`���ϓ��&,}�6�_0�X	T
���!�_*�@2���/%����@��������2i�Z	�1�����ҥֻ�=��&Y
s[��'�w�Y/���K�mf��|�(*���l9R!��@Zz���iS�"�~^�=���c��R1��SV�,4�F5ON��������*4<�T�<�����܄�xt6A��
WΜuܞO�6ܜT��T�;��^yH]�6Q����u��[��8�حaOe�f��c� ����:b?�� �Z�8_�2+A갯����(�0W�T��ㅂ?��N�P%�x᰷��	I�c?��鈫J#j �+t"���G�1sLF��U�*w
����2��j=�??-�y�y�7�w@x�~sB~�oU;k�5'tX�;B~>焤O�J)\[����N��C"T�p\�Y�^V��� ��0S7R~.L�k@hĩh��#+e�,�zo-9�H����m�c�Ё+^���0G��2�Nt����{[���x��!a���b2�.�%b�*��b��%aKA*)UF��;<R�Y�P� �-�} ��������_W�tF&��Q�.x��hq�7q�\��6̭�ݹK���<$����=*c�t�s�w[��w�[�3�՝�|T,��U�Ã����z���A�f ��C�"�/	��I�7児Ɍ%�H4~ B���U=!Sv�>�*Z��'��������{�� KbHK ���uJo�Ql��'ъ��n��t>����e������w��,qs��L�aͫek�r�hBbc�A߹U�C`������Rq;�@��(�
�\�-��(A��A֝�G�0��٘'�%v6�)��:H.��K�G�ڦ�o�.�C���G�N�:[MT��E�~T���t��ŵ+ܱ�|�:_%Ҵ^�������"�=0&츀JV=�)�V�T�u�p��6+m�0����(?�L%����2(ଷ(M �ȏ(u��Vg���x�y�|��-���	��Th��M��ڦ2�\[��pAi��t��������۫���A`�y֋��@B�ExBG�=�=����`r�:�?��v�Kb��LA�#{e��s�N�!D�� 3M����]� �/$�|�Ě9�k3��1�q3����RZ; 1�<Y2]�3����a�~0�q�U�ŧ誆�$�7���bw�l��]�jc�ow�����j��ZU�)��v��������;z�ʤ7�4��^H��U�Ւ��4��m�,f��h��ҋ�q�@��l��T�ִ��=>�ܕ_���*xX�ÆP�.�