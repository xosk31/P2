XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��CH�D<��/;�\x:��~FUs_����0�B�d�^��b0�B��jla���Y9"Z�܉y�cI�+����b���$�A���-)�ɊV��GTي]Z!t��g7D��.O.�z�?-H����R�(>L`I�E��I�����S��᝞�<���8�X��>�C���o�2!��Ķ�$xM9f�}��Ә԰z.O��@ �tG�O���;m,y���U7�n�\~�a�`ZK�7�}�>�ꎌՖ��8�a������8�H�
+k�����R&�����6���ī�XEL�N�u�OM�ğ�����3]1̆!��{t����u3��f���M���Mם��v�?C�ؼJ�>W<o �j�x���p�"��i��Lso\�m
p�fv�?H��'Q���-�$S�\o����
��!ȥ!�l:����
S�i&�$���_��A�������k��w�~���d
��/_;�p�d�cm�=�^)�/��]�\��8�O�Fh���_-���K���N���	sq�\��.��0�y�$�QwË2 ���dK{����C&N�����_���$Jf�p�p���b�)UN���Z��+����&�'����P���5ڂV3���r�4ܷ���Q'nt�'�����Y����4���z{��tq0ː��(PM0�O�CR�W�<�0�)��I����ݽ,��y���"������8ap\f��p�����K���C�B��4�ev�r�����XlxVHYEB    7744    1780�n�f3l��ˑJ~*���1�%yt-�h
_&�{)���Z&�Ƣ^Q(�L��*W�������ٙ�[�`��m�)7�D�^�������d�:}���1��B��=���]�v���َ���U^��*k�a�E�=���fhZT�Ʊ�Yɚ9�aoP"� ��A�lif!�Ȕu�L�V��V
��N�]���< f�(d�"�#�Yq��R=�hܛ8���(u��)	�(���u���Yut�
��+_��x~= ޒVNG��ü����1�����
6��ryAV>��l2��Ѭ0�`V�.�g�K��fXG�΁�SD�pXH,x$ac:�q�|��I	Xfn���}�������H�\�8DgD�2*��j��-,��,��.1=�x�#�T㾉��1)��䀘W���l��%�?e�rF:N~6n%9����.�e߅ސS���qc���� �M)�G�S�V8"u���^b�?}b��0�����EI�j��
�������a<�cR����-�w�Z�Hɂ��ȶ�V}ܛ7Z��Ubc#d���f��W}�Xu��!޳_n��M�#<�LZ��g����Gב`�+эB^�Ӧ�ښQ~%�.���;�=�@���a��pF��b`^�"�յV|�6�5�j���5N��M��Z��|4�"�g�2�|��~:�8�<N�2I���g��$��Ow�����ŨgdV�)�ĉ#��ٔ�
I�9 ��2 �^�4j��-U)�j:�t���b��L�Uq�Ą�/�P�֘>B�����Wɥ��r��X>�a{aT+����R�0& j_]�� �5Dy�V���)%���aO�j�@�}`K��į�y�"<K�}�"w
e�Ʌwֻ��.��$��Hz�R������ܵ�� "�Y�p��?A��aF$g��Q�m��K|�PYw�MStL^��MP�_���ͳ�Gu}�|i`�؈�xՙ�����(+@ ;���VNKB;ʘ�$�����@�Ĳ��T��祩$���P%Z^��u���8|[�������*�.����_|��f�W��R�}	���9f�<u��ܽF�4�"〾ʄ�q{�pKЩ0�������LqX�|#�k�rǵ�%s����(-$��)��T�R�0�&�f屪���O~�؜0����nY�ĭ(���f�d�� ~�9�W4��^Ѿ�v~$Q��wٛ�d�ΌN�:1(tW���Ȇ���9rY��g׫�h�ۭM� ��^�C����L<s��J_�Z�)�b�`~��G[�Fy�;��5�ʈߤ��,�!��WQ�@��P.��b������4.ۜB�6b�X����)���?�����c��M��:iă�r���&�k���{ r\F�H���ӵ)�z�E�
/��,	���R�	��ʾ'A �ň9��!:�a慅X���*AsFlR��U{����n�K*�~aK5�ϽAH���%~ql��+E<�b~�MPi��go*���8���]0�|"��j�{T @�L����g���oS�V��8�x_V��Hf�^Ј�ҟd'j0���5�\}�l�j"|_x��1#��a��V�_��
[>�`�M����`���gC|�4.�EH(����l��}��F�K�v��w)�*�u7+|��Ds�R�BRb�0@��[���������~"����)��3̐��Q(ś�Ȣ�/�}��zm$��c ��8lx�������{$��J��ҙ�"����;=�����-�&��՘v�>;'�ʲ
��[=��G���M���\s���Ⱦh�ץ�ɉo���fLa�4������,�g�{��v开�G�j">�bj0ƦA|���������YS�{y��4�A��'U�`k�8x����D���9����}}�E&�|+���T�����M
\W�im��ɝ`��E�G�+K��1��L[9��NR�ט������ٶ����G�8�F)�+�J�$���d���i ���YHQ����@y`Wu���{&�&z�f�Sœ�`��i�YS0�' $�걏c�)P�A�[���w^���F�iܩ+������O)8��%��T�!�c��axf�ٶ< �\y`��Z�<C�Z���3 Iy}i�|{�E�%!ީ�N?x�w�Y]3A�H̡H�Ix�]�E����k!��"�K}3�I�����<�R��L��)uRD'�Vg�ʌ� v�z%q��ǆ��k�����)��x�o���iN��,gIq��ʏ������#� _��4���W���6�đP���@��Sg�ix	�3�Ȓ��+��\�֑�D��2K���>aL g��[��<��n��[ȿ-z����re���i���&,�s�Lh���{n">s���5j��K�ǡ.2���ٕ04|w��{&Q.�s7�!%,��N+�նj@�c�N��%��yn�"���on��l;�Q���,�����Vʷ�Y2�|F��A��"��6���u��q#&���.��a��=�z|�]���$9�C9�(6ͮ��"b��h��FEJ�i��>"���蛯�t�~{۹��a1B�k,jۙ,^�f�z�|?uƤu�q��a�a( ����_'����3)�|8�-����xS��ߙ�}�lx#�a��bKƲ�����W�i����n�b�^e@!�����{"�r'�X\���	T�"|�&>�$������gӠ4nIg�����u��U1��o_�eFɻ���a�p1��I8��11i�����,�R�n�ewv"��ضQU��RKl�>Ka5����bA�@���{aP��B2�,���@Į��;��+����p��1@��eIN�;WX}�+?����T�d�Rmtm��[����NT����s����9�(3�Dt��� {,���5N!�.����^&m�4~��ּ޶��Lr@��AOR��xXB���u�#��U����jE�����k�a�"�Ұl	��g�rl1�|$��n�����u�fۘ�%d{*�K�O)�&`��M_� �*�6�9�Iid�00�'~���@Kr��z�����_�[�'�v�ɂ�,�~/Q`#I&��o�HZ+8�J����#܎�?E�T��Dn�xB"��tWr�~��ND;�>�1hC5<�&��6�}��+��x�0aoMk�G�Z�Zi�6L1 }��#T��xq����+-�d�����G'��@�?*U�8xAϕ줁\�oݹ���q���cΩ�ͩ�?��(<b{ey�>���_���b� �%R��޽P|�\5h̗w������/d>�Q�����?W�8��h��O����6ޔ�	�qH)u(5�k��5��bAT����S�ߡ;!j��c���FF���E�����j��j����lydj��Q8�$�CQ���kІ+vfܘ,��:y&��䂭�����ѷu�&���G<vԄ0sSnG��G/%���!�#� �9(qiLO[��l�t� ^+�ᯉ�E�Ì.�>(I,�(j�E�>������e��B1�dt ��$S�v�����e�=/�Z��Ｅu����W���Xit�7�J��+���mN���1kY�!S	9"�8UR�6��]_�Tm�G��b�,��ʋ�rK^
W��Ԕ��?���<a�ܼ���'���C����C0�]�>��>l.�D�%�����̻��~�O�S���8�V`��^�iM� ���q0_p05m��hY���t��16ݠ���a��L�w�g��~rJ��7�Y_�:�0׃�=D�ѭ|>LP%i��;J��-�b)�.�]�n�c�ZW=u�ޔ�l��]Ǩ�P�nk�c�N
����-�x�fy\��)HK��A20�zq��9�\ly��ڿ��^�|��G1�@�:���&��0�Ҕ�b NF&�~j��v!2��C
Ŭ&Rs��&��/���B��-�}�[t�� �����2iĨb�+�wSZ����v �)@��+�����M��B�OP��a�ɡsV(��%�o��HF����/�T_�
�E�rc~�!_	�p�����K:Փ�GV6h�8JZn�8?P
):Iց���p���V
^)'3�@0�|{���d��K�MVӘS5���'�y��$��3��H��x%WD���6��Q������+��uԖ%No�׮���  ��WBS>��O�ܾ�m�ք#˰���,!�*��q��OJ�P���Ē��������{�4OB�ƳN���)A�������:�;�6���/�{�s1y��;��5��D*��~�Q'm$��3�k���2������ғ�,�����&KC�	�J5{�R�9b��1
�؃�{%��8�@٦���]�CE-��Ɯ�Hޞ�g�&�h��
�+K�J�n,p���Y<:�֩��\�� z5�l�Ҵy0�E!1�P���4�N1�i��ց�����@�Z����������m���|���3Q���~.��X��E��=Y����c����n�r��]�{�n�v*�ՋP��S)~ ��N�"?F�ش����O9�O�F��k���j��35����K���դ#��8�d�W`�M-�a�Cٵ����-O���]?c��G�j��E)��d�cBX�%�QH�X��{�l�?˅�%�.�R}I��u����i�� ��,&3��c�yٸ�F���Kk�%@��5M��v?u�c�:_ó���T�Qz��9x#�yC�x�-�z���=�rG���Zb�w1�]���ٙLLx�\3���J��i�6
6N}��al�{6���R�r1���C,AU�Y���\>��U�e����S�p�	X�?��o��t���n�mdΣB��[�9�m���t�{e���	�"s�6�B�gÜe�P��䖽���.�+@x)���8�o4�Y49&���z�L�l�0*~m�Q�B"U@�g�P���ʜT/�EhR�hX������ґ����$��Y#������l��z�-�+��`"�?0���6�#�OJ���1��t>��?��e�D_�����#�"eEr��i>��~����M5%yϝ_�YCj�V	���B�����0�.�r��(�7�+��]ﱜ�Y��#���1P�tK���V��W�Z�1ǌ  ��Wdy�k,JVІ`O�N�gK����ϔ���9���x �>��Q���)��ɴ-�Y�Sĩ`�@��dވm(�ۖW���g�/�u��M���VW�5�'(�C��V._�b�Q��S�ʫ�EA���y5�A�Js���}$F�CV[�\�'jԵ������sI���ķ�0_����x���y���Gt
� ��B���ݪ<E�n�@ ,�߈�=\�>F��Y�#�]���Nϋ�eTv
��nc}g
za��I�3?��3��/(��R{w�h���^��f ��WSDO��B��R��f�m�cb�t�`7VyHEN�C�欢��ٚF|�O�Dju��u�~M��C���;���Юf�4k�A�L��,.��9ǘ8}M�v�0x�A$d���a��v7��<\BR�#�2W�_��V�3. Y��^�؋x	<1�cTu�3�I�H1D����z�qt���5x�=QW�<���j~Λqh!+oOY��D�nΙ��<n��_46^�&���#��.��*?��Twھ��ĕ�j+s���D_8m����*��]]si2�nG���T����4 �8��l��䳐�q�wU;�����{��N �����XxB �ˎv�KM���Ҟ��`�.�!ٚ���M ����gC��x4�[��0�g��ƣ��+�,�	%���L8�l!Dn�����C݆~W�����a��?m���oR�^�~�b�
ʣꦝ<?{7 ��#����e��`)�s���Eˬ�[+�m��d�@��