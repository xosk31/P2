XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��PF��n��{��^L��"spV�e�T�N:�&b�E�g��!:���#_�(��M����C*j���W�G���􇕬�� �Rd�}lGe�H!�*�j����v�ޘ� ��0?��_`���� ��Na��trA�=I�,b���nŐ8ҕ����1F`&�8XdEvJ:n�QV
��w�oY�1�߰J���"r�2�Zc�]�+9��l�����y�7�G7i"�F�[�/9����&�.
�(�#݅b��gҜ�)(?�%�X�[�ܭ��O�u$�B�����r2!�^�ܰ��s���	PЄ̔%��?>���x���0�wS� B�	=������/��3?DN�f���Z5H@U��yf�Ԝ�֝�a	ۛ_+���p~��tAE��1�9d�l����X��vMG(�)mn�Yok��Gwb]��e���8�:�B=%�1��M	T@}R94��T����h#)T�,��E��Է�_WW���g[�7�Z��Gm����y�k�oC��6J=< �QN?���ǃ��״�K�}�ǅL�aT0�d̍�Q�]wN�P��! \�\a+�D�u�T��;I����������<�˰ �O��ho��Bf�k������NX=��K���l�5�7�#���Ǉl�9��'�]�&�� �B��u	&�[��Q(o����y�Q-I��f�?��i&�����a/T���x6�g���~%?􋃼��������w��:W����o�'����Ք��x����z�XlxVHYEB    302e     c70
yh����T���	'�$��aN�"�{�'�ə7�9F��t+�������$b�`���2A�h�g�@t����\�u��<�<Ά�w�<��++bq��ְ�ke��Z4�e�L?G�nz�dQ�3����\{�+CE{Q�N��&�F�,�������1�������؝�&P��(\g�|��A�`���kQm)�N���<
Y}먃����^v1<�����[-쎴�瀢�"��%��:8���1�I�0��(<}pmv�]	e��^_7�>vtt�}�>��tdE����&��p���7d�wgm���s\��Q�G|�3<�L5�F
o��{3��e�w�B�K6�U��� �h�'���a��3\ch����B���霊$��ύ3��R-@����:0u�8��\z�����+'	���f8#�NL��2&��Nr���ZT�h���m?a��tFʫ|���Ȟ����J2�8mg@p��]'T���T��Aj�/�W�+�C�fH��Ҥk�u\�����e@-[�Y��kG��D����?+,�%�-[][^?&&�3�<f��O"l�w𜳧�L�S`v�g�0	4��5��fA�o��������-O�]����2f1q�3���=>8[g*BD��h}��,kF�Au��,>��p��2|�:��8D�$	ܲXT-�Ơf�Œ��;�8�f�0� /0���$o��4<�����V���G���^H��>��M��U�5m�@��)Cͮ}4D�ljʢ�]d���_�B���1��$�H]��W��n�81��vυNѧ�x�,�d����k.e��_�2X1�.W;}��x��fl�n@s�hX@b�����04��f��-T� o,����O�k�vnl�+w�H	\�)v=_vV�*r���k�V�WY��A1�����_���7���T��NaTKe䇫�����`��|híY��P��"ܽ]�m@���V�Lĝ�rMP�m^0�_���G�i̔a)�Hm�d�9�"�<��t����i�<��=)�8���U8�VM�Wĺ�:O��$��h���1��;q�a���Ѐ�*@6��E��#b���*�@������hY�<t�9Z���=�%\�X�ڂZ��80�2��f�F�b����y"�ە��c�t��<��]_0U�x�+4�n8;~?�����}��B{8 0o(��7�[-cnz4J��8��o�f���3O\'����i�<H������fm�6m'(A�]Pv�.�>�_��w_<���v�2��зe�ұU�T��Z�����`�"$;��< R�w��j���M��PK�e�A�w�zëW�oZ��,H�U�]���%K��W��pEHN�Be:g��^�ʻ�A�b�Ց�]�rMށ���ym��E���H�`*Q��l�~e����ۈ.��8����t��+���g<:hA�f-�����ǳX!d�%���Z��_�i;�/�
鷎t
�L=���'���C�`S�����Qu��&w0M�5"�_���(�k\����Gط���y�䎔��C��4�?"���|��������gw<�Ќ�C�P�	�,׎��~����
�e��y�(��ȟRyH~�-,B��W�� 4�e,?ܐJe޸M���`mEg/��n����f\�>>�lt�q~��h�U�DPH�H��?��5�;�O�0�}��P����F�����p��0͵��]�^�=��]���E&��L�k�m�[Zy ��g�J�CUWV	�`��j��m�.K���5��>���8�t#�q2ld��FH����_�[�1�'�A���4�2�(��k_AF˟h�v����n�7���g|b���5x��.~6F�e'�D�`���MEe�m_=�{2C)"a�C�
%&Q��|���sp׳��=`S^��dvVP���L1�@�+sg)�y�a-.!y{NY&&L�t�u��(�B�Q�_�9���)۷p�n~%w���g4�1`7Aʇ�|������r*I�\�LKy��d��kbv�i�7��H�S�D��~�CAmG��2$oRlo2\�?�Fvv;l�h�Z܅ ��!���3��B��/>$�����¢_Nޥ]�ʝAD�Q6���4cx��[��T�Uw�ۗK]��Z<����DV'fp�jK��iI�]���o.�d°$��T,�W�Trڅ�6�����N?s5����a!)h4
��X3��M~��8�&<�J�4��Kb���҅�H�ta� wS���8[0����!����lye��q]|w��]�ޒMw��lbt��rI4@�����B��J���l��/Zj��b��2��
���SK�]��:�Ω�d��c�����JG��3C?l�w��38��*����j1�!F��<kX�[��zMm=����U�ъ%���&yژ�����k���%����i�óp�����trUJ6ۿT�ݠ8�'�����b �N-nIbm���%���y#�{��/O\�Z��Z~�U��Qiw�Ӌ��Ly�]�A�db���<v��ؗ8��B��^�U��'sp�??�Tb&�k�L����/� �R�M:9xE��t�9�ǁ�_yF�S�]BT3�&�V���L�,%�Mc8i������L�irWL�P8a�%�e�/����ާ<�����D�Ni!5�>U� #�#����̀�L��Sy_��&��1꘵w������4f��7�:�/�sڞE�h�x���.�&�2�a�mz��?L�s �w��K'�y:�26�r��ؕ$p�g���c���)@�ި.�*j%�요 ��>@�{9������0�/���l�"�6����hX��G|�B~��w6�庞�$f��K�Ӻ���,�w��p%�8��
�Q�]��w�Q�1l{T�~g�K��;L[o'0���:�.��@s��M���������.삿D�W��2�j�)Э3��`�<x� ��(g�ϝ�S�p"��>H�!2h��v�y�� ��'��a?�/3Ԇ^t�L�d���~� �g)�wm�T�ˏ�A����J`�v���ND#��|Z�3uv^7�(��>Ρ(��Z��}�^~��&�O�O$�{dn���?���u��~����@�j����e��Z��"�S�