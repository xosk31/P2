XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��\�����eS����Z�����q�jm��',m��h�:���Ҫ���vD�fc�TH��cD�T�:�C\ _�O�*ފ���c����溗���%���} �(�O�,�_j&�<�� �
yҺ�ښ,-ܻi���%���I�@��B_�7��Ϥ���o��.~�8	��=%D��ʺr+.g<c�X�O+��(҄�5�����:YW
��;�/��\G)X� �IF0�A��'p�`�?�O�e�Ɨ�-ca/8�߇7G�S��^�Ċ��w��4���"/����a9LO�P�!cvR����ɝپ����@�o�z0��ýx�>P��m�x����h sV����cV-���z-�Hm�v��j�ڽgڍ0����Z� ^� 2����T�A*��PS�^�
����@���r��X�������1�g���n�(�g������}uP!ءs'�
e^��!�Q��9u̧�Z{��9���9���׷�f.�+���2(�-Ŀ���Dj�Uٝk�����Z�-GlS�!zgr���f�Ų������x1\-P���ӎ��m���a����p���/À�U�i�-D�
�8s�ե�!�֪xF�1�'��y�Z4L��˫������J�:/�Nڮ�����u��64ӭ�	������CB[�/	9U����~�)7h���\ߨ�m��}f6��#Q;�n��ʹ6��vP�h4���F��_�Wa����zTIj׳E.�����A����O�!��r��XlxVHYEB    4089     e40<Z��~X|yz8@�EQ��^c	^,ʢ_@d�9]4�Kr��t���.�6�/5�-��:r���#1U\r{R+;�`OF�G���ݳ��𼬓�gy'c�T_WkϠ/�'�9~tT����շ
A�V�<~�WǊ?{N������XPl��G����	��@*�DK��_'8C����K���x�o��5$ͪF/0�h�޵T���^��~��Z�@����n�5�7N�W~Pq"΁eN�P%�oa�Q���V�r �K�]��~T1�'o/>T�,.��> ���������z��]e,���L�m�@1`��+���wR�f���V��4�Na*(D�1��K���D�j�&?Qgpi�N�Æ��dHZ\�Ogzxߔρ�D�ʞ�A��x)A!|Բ��Qy�o����T`���"V�"�;��(�G��d�TF�K1Ʀ+8��S���������*��R B�|�; ƻP�vL�r�1L]]�Im�Q]SNA�9�m'ᤳ�ă#��{"��ꌥRH(��)X2V��Q�ou�"V��y���u֙�������N!{��̇�����oX1�M��{K=.���o��a���<��:����ʊ��y��Esw�D�������ʷ�O�с��  Z9QCl�L���l;Ŧ>C�QN��LA�	u����o�*wr���Tej"5@l*�k侉"6� ucc@�e��aIL����oԚ�Ҵ��Q�d�W�5��\?���y�
J8f� �ǉ�
��I�\q�������*�ԩ{�a�O)��j����LB�R�$�M�ᐗ���Z��`�Nv�������8�P�&%��Ddؘ���yu��z�i	���mdu	�Xngr;/Sy�pLz��Ȝklժ�b��te�+��8�_��|���:*��U�#'o��� ���xV�`Q��/�҅����g,�܌���4���]�)	S��i�tz��A��0F��N�^��-�8��kK$��,�Cx��ʞ��^�/S3�+Hdg�a~���$��I�*>��΃1hx��H'�����dkQ��Apt}�EEv,����̱�~E�}|�X�ļ^���'�㝶��s7�^b����ʰ4U�r��˻�Ʃ*p���P8����C Xpw$ �ْ3�=�l�Iy �.R����$>�k���Y�3�5g��Ǯ)	=\qW#:J�\_)%�h�vk�pz��o���功>�"F�7�Iʆ �M��/�W�'����K*��À��e��@��|<1�r@Q���#�<���7�n&b���"ɐ$�����)�+#2Ne���%����5���e�z_���%�����`���߬�ó=���F���� �P����s��� ��E� �)�3��A��v��#u��5븥MA���2x%ʴ�޺��c؟EÉ�a��l,Y�bH�g?:��m3�~�q4K�A?�p{��i��r�!Ն���Xlq8�4����z���g��,`�R2�h�|.�@�~��KQ������Ѕ=j��U�ߚ�E���.ˬ��+X�KY���n98��XI��%�����M@	�h��p���t6G�u8��j:�/,�W[6��������L��4�G
v$�����uy��	J��ЎE�>?��M�� �ɦ�2\��9MJ�v���U��,�AQE+T|��`�O��2u� �"�u�[����>�	|쇻��gx;�FJ���p�?PlD Ȏ�V��dv^��f�7��K���q|�$�.r����N0�U#���\�R�s����1AɛK&�_�Jt��;J�Y�%��B�{��s&��_��,k+&:5�Y8(Y��ʘ���VެW�?��-ڛ����~p駶�)f
E��n��>��D��a^���^n08~�%t���^��U �[��Eƨ��F��7�JL�6�~*S�y	ă��s��d ��:��3��k��AdL`\������P� B��I� �r�'���5N&"�Ē�T
�C�^Q�{>ao�G�������i��~o���+_�T����7�{s>>�(�O&wdu�!�P0�R�-���ϻM��0��CC`MI���v�x�/5ib���}�E�KU�x�.y*�e��vB�)D�k�7����V�<�'��W�{��9Կ���������C�a*�X�F���n&�g��rJ%O`���Ey^=[읏o����9�J(�]���уϸ��c�֧�QDv|=-ޝ` �;�g~��wӒ��Gz��M�cH̗�Hk+FW�X"���̺RI��E�3��_�
9�\F��T�X={챎�7�x8���U�dO^O4�k�M^���O���eQY�lc�f������3����G6�`nO�譬V�5�b|����Z�̌:]��	���	EFxM����������{.�s�_�e�FC����IK�M�&�b���C��Y�=���ץ,^�M%�-�u<��f�w�~ȓ5��L�,�2D��IK9�I��y�#Wd+ԓ"�]�˖������OW=n�T��S*o0í�K�deZu��J�Yeu���^Ғ���v쎑|	��7�������.u�w�웽�k)��E"��Te�s>��J=��D�g�L�㾖�D���Z�c�?� �s/�QI|�6_:�
�^�$D���Y��j�ٯ_� wH�� !�\IJ�p]��m��6ن>Da��v�?���Y�O:�j&&�:Ӊ����z��/�WXD	�
�M�-�=P @����E�W���F�W0��k�j�c�����(]���ɵ�Zl���r..��t-�4���+�Q%�q�#`v��|��+��NX��[����~s���d%�Y<�#p	g��):+]Z���CZuU;}����c���!l��uP��k?۔S��uO2�S��_�>Ixv�"pĆ`@h����4�c�E65��Mn��K]�zY<7��H���;���#(|n ��:5���^��ƙ�7�he��^6O�Ut.QEuS��3h':���˜�"��	�Z#x���F��St5!��Ҹ��0�c�X�T.ڰxn�"���j�nz�YY������1X[��9�V�+��?Y��-ak=@��W�I��#�6Mu�C"QF{�A�{��d�V���MvDT�o�,����Ak(���E�B�2�$�EF1ʏY��Et�wB��n��
��Щ���
���u�/q��<v���)7V�웁�υ5�b�w�{�qKj�9Ƀ��a�U&9��"G���A�2x�S ���C�����|e1v���"��]yعP*y���(�w@*�M�%$з��[��B/ϕ�s�8���d�u�B��w�i�T
��� � PE%��>?�-k�n;��I��?P����m�h����0�,/3.^�������Bw��1��Q�[�3��Лk��,{��c�wh�;[b$��z,�+�;js]	e@�3�C�e�s�+��J�$��M�ġز�DH�q݈�5�gV��:���i��^%�u���*i'��w�&Y.n��ǜ�r~��w :ʳNM�4g�rC� �T�bU�]l�S��Ed�̹�s�'