XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����9����|j�I��s� �?͜��I:9�S1L�n��Ee�;<q�{��ܷ��W8���'��j�=��+D�z��v�+l[�M����9�Nl�	�S�����eXF�o�e1H�b���uevty]�K��F�¤	��Պ�1Rjg�I�/rp}�dKNA��1��5��4q;2[~�7�)v�`�cYa%����:����w�g����ʐ�U]-ʍzf����n�:�J���I�N{|�h�D�#���M���¼q|�T4��2��q�2:����#��o0��1K/���&��y�Y�5�(���K�(c;}%+� 6�*21Yre��yWlɽ�<�x=PՑu7@���hRc7�q��U��m^)������W�?��r�E�9�������+>�����ѿ��� �e�Cxw���J� *q�V�*��(=2��~��j�}�%��X����b���q��;}��	u�GRrp���)a���<��ҏrw:� �\9߀9�1[m���6��/�΂B��yh&䈤�K>�ι����=��$���9�!�R�P��|���F��	7	X��fj
���%��Ђ���Z�ۜ��8�d&?�W�8E�9��WZ9�A�H���l���L^Be�r�[Z��?��H�.)����m+KyF7�ωW��pO���z�I�@��1�)n&�O���o���6�*�j�ss����6�ZZ�q���Q�b)@ ��9�~�%�P�� �*݂2!m��s�9V�y��(�XlxVHYEB    2dc6     ae0��C�@�	ȕ�k��>Qzc�����ա�.�����F�O+L �S�O��,�q��6�=5�������e�"��J�aG$x}���A�N�y,���ꡍ<㛆3Tg������э� ����
F	�~��/Lc��'��PA�Yze�ho������ϛ���r� �*�=o)�k�Ԗ�Ȥ!	�k��}���/�ą�:f�.���d'8�k4�^U�=-���#Ȓ��ѥ������*����<��hX_���}5)�$�p��A���ɆVs��lSe�8��q��t;4��)��b�a���X���.Ci���0_:���e�kA���h�=��U��1��9�3ē-D ���v��?<sEɡb�)�B�ܤSIPoao�0�� ��i���+�7��Y�Yq:�U��>��k`Wx�u�Z7�p4V�E�����8t(��G�Gd�'���|�� d>��ēoX������D�~�L��I�K�����az\������,)��_B����� p��ZD�|����SvBڙ��#�a�B�Q��������8u0�o�-7�ӂ,��{�	0�{d��q��o8e�)%}��.2�|����oU�-49#T��?*Κ�v}P�*U{�JP.��4.���=4  ���J��3�C1������nau4�1r;�ǉ�*I 82Au��ˢ�ZG\���y�_C�B7iO���d�S��*5#�Mc��q��Յ�����o5!l�r-mG�T�\�KOR?<��=����~�1r�<�L�J�Ƹ���i4�m��s8Qe3P��4�?[G�շbv^�_�k��a���˭e���w���m��hC��ugszg��nHG�nb���d���-i^��b#J�I:�cI�2�h*߄o��R��UU�,�d͎�_���V��D�4���%��5u��W�q�F�R��9e�MͥD��8��Ŝ�:r�\��IەC.�2#͟�<|{�Iŀ���c&��gߊ2�u` ���V�%�wv/�/{Ł�����S�PJ��q��L�U�]�G2[ئ�����4ٕdl�}�(��.��Ē���$!��I�u2N�J������g�տQ���<?��r����č(y�,�b�5��pa���|�˙x��\�W�]e�Ee��C������\��Z�ow�[���-LխR~#��Ifƒ��b�D����z��&
���.�L����@��������qĈ�P��o��!r$6���"//(�-�i4"������+��R^	m��z��,C?:R#F�1 ��uh��غ��J�~E�M)Y�*ۦ.$���@Cq�#���^����I&�|��;���V�
�]���ѽ� �,2��Gj�����
��hz�c�ƊD�R�VNQvL�����iEs���,�����5"�,���p _{�V�5Y�U��ώs[k�t؎�r��tݾ���� � /������F�!�4�r�� J���d�.'�9H��f�х�n����^qc`�u�BЁ�����C��x>����>�p,Z`%z�F%)cK�"���`yx���(��]�2޼C/Ӳ���|2��㬔�� ����x4��<i �M�����W嚗)�M�k��q��#bi�>6���*�v���1�ߚ�hi=KAn~ys��yq m�71�n�b.�M�9M�r��;&2���L�-�B��~�Ł��mI���p�ZG�"�8��f��H��qD��&����$�#c(;���R�.L�_䲔Ad�&Q�W��l|@�f4�g��hLEU�^hr(;����[�o��"[�FV.+�ѧ��]��l$���x2<"st�9>ro� ���Y�Qp�o���|�����nf���Յ�X��Dػ59�� B�������n*�i�W�[ͪ��Z��4,0�V��"������
s6_�6�`l�#fsgč���5��Zd�~�Rhk�u�ק��hŰ�sK��c��?�� ���j���-�C���GE�g�hp�"���k5�{T�<+���d���96�N��s��8KF��u�xC���ls'v� �����6�瑖�ǣ���)dBm�a�uهe�WX}����Л�|ҒoFf.C��<��g��7����QC���N�?�l�J��J�����Y�"�zX~���32����|��w����B���Y�q�R�۝�a��ݜɕ\���|�F����/���D��iP����+�r�׼"
B=��UPh8�^�m_��s�8"��=��$9�x�,�V���)޼�EAI��d������*�$M�:�~�m.{���6�o�̧��T������{է����q��;�g/����c��t+�� s#4�4?ƥPk���>�*��=��K��aѧ���e��������:e��x{�ye#HK�"Np#</�IJ"�0��W�B�����~���/���3��SwJ����L��nh���W��\r?9A��^��4�~�A)����w FMfl��O�N�d��Z_i��aA6Ji��j����\r�Jc��G�E�FZժ�Mf��\�"|�X5"�0y��z+�i�0c����|"�">�%-���E����M���P�ˈ����#�!w�Dm��50�3�-�:�������d�s��\�>��uSQ�/+]���
*t�@�l�PG�cǢRҭ��!5D�Q��a'K�ȋ}[�����<0��~���Vu�~