XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��9D��s���2fm��U1W�*���wl���ݝ�ks��ޣ��c��X>�6u��B����J�������M:��k=�s�����?R �j�
}K`�@�3��|T�Rp���?-9��ѓ\��$ ���}:�Sǭ�s�h3�z~�`�%C��O֘��>xCq[�.ⵌ�P$Q}L�G��7X��(�s�>�e8g/XvC��8�/B���JbSܙo��
{���(�J�FZ�e����A���a<J����
����hs��0I��w���G��~��N�]��vn:٥�|h���R�#���7�ݡZR�๱o��;��S��*Rѡ��j!���5t@�dKk��'#��e�З�*ܒԉ�XpYo�5���4Wh�À�b�����);I�ϡ�B���D�}1S*]���� '��7���Z&�K�3��h�֭�韗����b;NO���l���H\�%�_t�W3�<��9v�w���"�����iH>�ߊ����-�+���@� ���g�li�GӶ��3ud�����8j9+�0��tX\}��(x�W� ��q	�sfA��K�q���wo(�q�ٱ"�����Õ|4Dwb8��%U��L-���Q|��V�/��F�/�L��c����tx8����{���!�������⎥�:�f��K�9�G]�d��&�WqA�y��)+0*��TfӃG�&��s��(siY��=���y�>[Uuʧ����[��D�R��XlxVHYEB    9de1    1670Yŷ��_���I�/�U����w�Feՙ?~'��-)SLfS�u�	�.����'?;� 0R���&�+��妴���pI	u�����p�fC���65)�fh}�A�����m�ۂߵ����H�b���\�Q�t�ɤa���*�im-��=���\�t�[��� ��%�]F����WMVT/�C/�}~�}��O�,�3��@���������$J�6�@��OH�T�7>��'0����L�;=w�T 6^�ɘ_���O����4���!�4�������s��x
�|_|�kv�2R.$��hlk�(���hdT�BS��c�L�����!�ǻ�?�Q�b�૳F�w{�H�(�I�y"�4���9�kTp����R�䨢�G��g�N���?�6 zxb[2J�	�o�t�I`�=,�	��@w<�)o������Q�ê�E߰ON zN㒅���H$�M�����vw�z��ӵq���̯�"�(F9�x"�u�C�)��:(�M�W~�V����w��m�����R��6��"ؖ7�4��`_���������0������?�����iq�F��`9:
��aM����e��t��"�3�f�2M�ؠq�0cc��${�r��1!@�@f!�Z��^�������ϭR�F�YC炷.��
�]Zgh�7����_y�aF7�k����T�-��W�M0��g���@h�
a�$���`�æ��Q.(1��괻�VsI���D I*�$~�mҎ{�����*��S��4j�zв�׸�Dz�y@%�^�S�D�>+�F�O6L���Jk��j) 8���!۶�{��p�Ћ@�w�Zft�׃h�����n�gL��3%ROKP��B�^˘�������@��x�C��݀��L��(�����W��#��!�.�`�A�a��g (E�sդ6P&����de���\Ґi�rƳMZ�:XQl�_��mf-4L�%V�vs3nV�2&���Q! k�ߌ�!�=~��A#��eM� �v�J�i���1���U��X�,���6�����	썕���6sp��f�S�+�nVϫ�?v�~���dq���# KҊ�"� ϓ�ƪ��� ��?��hF�@�v�Ļ/AjV0v�.�~ӓ+�(hUa���.��S�"�ڤX^F������U9l�U�����I�uR����'op�8�g����Н"��5�Z�N��C!|ڶ����!�R�:y����� ��\L��X�R��\1z�l�Y5��	_0? ��͵�g�I)���e��,,���%�K\�wE,Y��Nv��kEub�ʨ�V� T>c{��\�V��x"L�'�/�t"�ಱ��zD��[��,P�'^�xkcF��4.q�8����2i�[_M�V�6��F�ۓn��V���Y:>�y���s>���C�ri������3���Id�M�����i8��?��,瓌8s�K�3�e�E�=�lUY#(G0�z΍�r<P��}f��M.<�^�]���d��E�G�k̏[����.�F�wW�\:\��m<qR�SX딹���rZk|�_�r�x���V4��Ltw�Y��O*�m�8�\TYR�uXWшr�4�fD�w��`:��-:Q=z��8��f/�
�^b���`�} z�֐R��jOq
�ݭ	��ۓ�C�6!$ON{-���]�39Lߐ ��뉈vX��M�4ETD"��w|׈C��*(ci�<�@�P���Q~j��A�إ�J��1J�#��h��ZO����%Yo������fi���S;Qz�x�d<3��2ۿt*�1�YpY1;'�H\��G����]H�w����@���D��2�3*_��*�%�Ql+8�3�c���^;9�h���L^�7@Ґ�T�U���{�Vm�迟�3d��xK�~����o�\}F#sB��ܲ%ǁ�q'�:���y�ô�|v!���et]nIQ�r��d��'|}�V-u�r7��K�$*����Mfn�~����q �D�/�;��4i*$H� :���ߣś&��L�j�0���$����l�������1��"�=��d2�"z+�\�Z��c����}7���L	H��F_2!�L�E�tb��8��䅜��4���"`V��MJ�Xy�9/�����s9Z-�EbN͌��S�>�j�_!� ��g�Z��V���-`0β��1�;Z,��Ϸ7?lCsY���~̢9�	o���1��f��o"^�?��o�~��>�b����J���so���f��x�ܖC��ӆ\�씮�K�ڸ�£�i�:���# Jvxzmkok?���H�-�ؿ�Q��|��\;��?ᰍ�'{�������N]��^�C�� �9,4ƈ��JK�zQJJ��-���N�9G�v��m���Ɠ�Hy�9��&_7>W5�|�T�����������t�Á��rN�vK�.>���l� ЍN���Ψ�%x�"FZ0�px͏N�n�������I
t��A*����	G���<���d�C���ŕ3�j�����5������ߖ���`�nYW�-��/�����۬��	�J��w'�DՈ@�[|h���g?YH�$NɭUfv�y�����3��u�[����8 ����|/yc��� �^��nF��N�wԺ0_��>�>09���V%�����-���6����&��ч��r>�C>��rǚ}���=~ޠ; ���zy�?��\���m����U�x��v�=�˥%oXn �4Q�袞q��n{���d�"��j�X�p��4s���M�-�A�2{
���=�v�+�.�DdD�h&Ɂ�:=s��1:K��Dx$�et`�:�$�lX��#0��x{�-���2����Y��E�]�4���*
r���~���� ��BX�u�v��!;��a��-��<~}qy�����^�v	R�
Q��PE㠐�@t.���!en�ߗ�, �(rxVH.?=8hl+��{��I��Tw�MCh�A��it/$�a�G����n����F���� �)��[��Sʭ>�/����?�l�%����3*gº1���(�Tߴ�τ�ܡx������P�!�<d#��#;eL�fM��{=��j���М���ކ��
�$�bm<�h���A�*��S�n(�����PB��ф�]�r��w9�/�-�m
K�J�o�o�u�H[�y����HJK�����2LM[��]}ɶ{KwBr����Qm	!�U�5��?��dJ�,`������Mt�� �oy�8�ï*���g�{�|��t�~�W�k���){�L�X���w^/b�q�����M"m����]PT@�l�'Lʀ�UQ���z3�Q�"�ux7��K ]�Y�X�(˲�Q����[4�%B�j"�#��b�9e�_fm&͵��ت�'S��ƏW��`�����A��n�6/�K�0=�4�WlPZl�QP�V��Mă�|��Y��������7s@Y�w��`�'Xq;F�����uq3.��������a}74�v���!��?)RV]B��C(�m[���᧗!�?A0|Z ��u��/����{o��Y�kLdcn�sq2��ݴ��N��!S���+����<���I9Zi�0�>�]���\�Ϸ5;;�öWcu���T	��x��XT����5I~ /�q��l��$pQ�*i��K� A�ik�h0]��R�Y3�$[��VL�&q,Tj��[p2�>4��z�Ћ��Za��� ��"������0�Sk5�)t��@�3"��g
יb��q����L�貤�H�Qbq�8����3���p��(��+B���m��J}o�$;��|�$�n���O(Df�"�$\�����([��$%L�z�7�C��B�!�2	�/�V/� �e�B��і2��G���uy�9s�y)��u������Qh����;�&@���������z����j�"q��zR�I��1A'��65D,�%�!����<0�k�����u��&�V���^+��'��(R΍<{B�|<�z�$wdڳÑ���1:�ov�D�f���!������HR4��x��4�0��y�B\l���Yү{��>G����-D�M�a��&]�$���}�b��;~@��l�Ͼ�$KTs=$9?pOj�ч��8E;m_��~�ǲ�ˠ*��o��=��݄^�娱���xJ~���ʈHs�M����s����U@1���|��Fp�UN���;l\�=�;Dk���1���E�`R�F;!e��F�@g�S&���;_��c�{z�.�r-��ǋ	�{d��̦����F�r!M���l$�{f�4y	�A�h����´1��(�W���ػ]��&e�-#�5���`�	���ߩy��'�͊�|c���!��kcͲ `��(�f"�&�R}�nH��I<��?�?vtԪ�(�4x�G%Rѡ��.�#of����c����V�u���&ۖ^���|��༮͵�k�N$T|g�rV�b�t$[�0:q��j��a]�_�lǂ�$p ��T�vȁ�L��!
�Ԅ��i�@}�E�x���$ܳw�����Bg�;�w�$y�i|���� b-��qE�3�-h˅�cZ��.%�����֮+�Q^پZ�(Ron]/_���.�|����`'(u^�v�x�0��'D}R���Z�E(h������_k��	�hΖ�X#(���'7	ˀi�H�����#r%kG=^�C�&��z���<x�I'�`9�@ջ�>bmy�0�4*��&l��*��uᓾa�� �:%ò4�7O��JI�8!�(e~K�K2���Z�\�G�p��l���Y6�5��K�#�h�8l�� ��m��(�w��Ts�t��S��Op`�$�lG{G��!�I�����y���S�R�yXF@��C���p�@�[�����)#�7NA��E�+U��9��|{�$j�ٶħ��3�ۏ��
4E��6��%B�EKk!`�'�8*bq]*�8�����!��աƒ��� `�r�?�-5s����=���:8���M��"�5��š�:	Y}�ً����$�ƿ%V�94A"�nj�=鐒b��� z1���[P�#a;��rs���'�ϝo> �F�@�����)�u��fq�\]͆�M�����@��XG
6o��YmO��l�[Q�}��W�3O��W�S�G	�7�"d
q��_XTK+�� �Xn8���e��~8�P�6�y.����z��)�O�9W|)P	��שb;��*�El2H�i㼦���v�瘱��U�V������4%<��V�R�8�ZKR �H<e�ǼF~�j���.@{�?m*���3�o����`����/�ǃs������S:.ݮ��4O`٢C��|����K6��M�
�A�@IG����Q�I����|"�` Y�I�'�����?�J�<�ʆ>enQjǰ$�܆��������EC�1TQ��Zqy��}iX@�vZ����G�񿊵5E3�4�9C5��͆��6���O?̠��3�|?'�<ڽ�E�A�[����#fWt�a��#oE[��Ԯ�S����܂�M����(�4L����+�^�3�������uc��h��`�p�X�����