XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����IYx����Y7{C�ȏL� �'��mq&�e�poZ��`��K�T q��s���5v�T��0��{�y���ߛ!k|.{�*\��+LrHT[phx�Ā`��@�*��t�F�аj�~��t�V���i(�����"��XJ���W����Z�4��M�� ����9k�C�oӑ���GX<>O~eA�@��6�'U��h"8*�1�n��ڑ�⹥��z��o������i\�����6�/q��ēt&Q	n�Uʍ��vy���u�Ưg;ձ�Ƴ-XO�����e�����u.�c�2\����j�}|I���BX��@U �p���3�m�ݭ��4�vX�tz�<N�E�� �<����Mڴm�r
%�����%�2ar����Z�T����ܗ��oA$s�`Jέ�e ��7�P�c&�"j)
N5NK��!���2�������7I�v�C3oC���xYc�x���;Y-"���(��lT'D�`njdL��b�Ok�sof�)h�eQe��_B�"�ڀ�VX�	��Or���8���r�/O�OX��\���X��[��n�8��4�v���(��޷��&�mV�q�W3�%�-���K�f��lu��]mIy����Q71U�)��m��17Z�\�:��\���w��rV��L�)��.EDWOSl��X���][n߷@��Η(��w�8`4w�|!�m� t�k�ێ����Lb'B��B�+^Y�;W�nPگ���`���wO�נ��5�TyXlxVHYEB    da14    2390Jb�~ÍC��	�f�+�PՊPQX����_�:W(r��8�o�_��?)UMU�!�a!1���N$�������qu/��ɿ�t������Y�m_����\�����Nu���O%���)��N��w�.ͭ�W�Nr�+|�f�(S��L�Tڥ%Q�T�>�5�Jgj����F0��T���{�L�a�B��F ���aC�K,j�A����Z&-��:�F��8wU�5�<���f���TW�		l�[����e��z? �"!�΄<����C8P��|��I��*�W��m���m���6�방�9�����n�#2��!Z�ݝ�*��� �&x]q媗�]V�h�l�z[��SV�D��`c�C�P�:Ȱ����ҙW:G ��֤����|����.��#_�(�Jk8��l̰GD�<=���0���S���D:���A(u&e��C��_vJ����A�{���B킋����,�T�D<C][R>T�0����9 ��G��X��)�2�B�{U
{����Ꙟ�7��l����I�����$Z������M�9�E�?X ��x�(��ߺ�Ħl�	��^���ꪱ��4[|�p��Ӛn]�ۉ�
�]|3�:�º���_3����n�W��?fG��Q�tR�xʹ8�?���;�*@���#�(]v��F�=h�S��/��ߒ_�{\��X��Ћ�j�*ç�}%|���9��w�'q������Ju�x��_Lg��M4�+\�%]�I�������Jܜ��Q�.�-�)�����٣��)1�f#g%���~V[B�/��)5�H7�]� � ����)ŀL#9�����2�75�J��q�r�G~��[U-\�G�ŀԬ���?�hw�%7�P\�����&D�+�˺�/����-,�V�X!���U�@T�,n��G3[��M�\���!���ޱ�;M&+mc��(�NH��[���_�B�{+�.��O0��ײ��
Wm<`��J�q�!��tp�X����$�BĜ���7���\���c���9�,�t���/sJ�߯+��_�3����Q�����)h�D�Cj��8�`�Z�ty96��Kb��-w<��ŠQ�/q��)�w��!0��m���Zyܥ�=�h��Q]��3�����{K���h�[�gO��3u��b=�#�N8c��Nm:_��L�Rx��Xs־<�91��o�`�u��1���\P�6b��;R��B��w��F4.��o|&��1����0��ļ2Z�P��xNB�P���*=�P�ӗ�`ވ��0�0[��v�Ȗo��o�y=�[�GF�WvO�����<[�����ӛ⏔���*���U�6Ġ����F+�}G4Vl�c��U�֤}���@�3>�~��/7l�g�B���z#l_d4��:�7����t�	����gr@�JUП]��m��������܇�D:dL�~���d��&DK�e����xC��ў] �ҿC�\q�̛d���_5���PQB��l�+�w-�P�N�����_־j����q�=��R���mR��2�E$w�D���-a��j�rǘe�z��P����WTȸ�?ަ�j�?�2u6�n�g1�%	��h��;5��c�H��_W�ܳ9Gӗ)�]`S�C���L��DF!��.�aq�C�p+g�O�u��]�q��4;F\���0e[	,e�F��>������J��k�bR����H{ːeurP(���Y�_�ۿ5}����ae��e�9��~�u�0�<��y?<���g)e�u�.��5��%:ڠ0+P���;�i��M�}y:!H
�DH������Ĉ�<�p&�<�	��>tݔp�\���Nݗ�@H9�\�s79�[x�U���߻	�{������۩���>�����e��ݦ�������}���9��|�a��xbe^o�{B�0���Nڗ0�����dڹ��뛙Qó�3%�H��
� ^���*�g��Lk���߆��zh��h�b�T�d�ttǥ���o1��+7�TԪ^P�U�b[֡Q����}��L����L�<����,�i�@��fAk�c�L"�3�1:�{�, �K���h�L̞���v��WbFZ}>�)a�Ɲ�Z[:��\�x�����?�c� �����W�.B���^+�3���,�5���3�1�oS�*�ԐTtp�;���	#�fB��6����e��=���':�����{�����~A%!��e��זR�z�T�'t#�gV p�L(��W�����5<�}�Y��]�r����̽f}��r�K��\��%OM�~����6ǌ�L�����1_d���ɡғ���������#���aj<�2j����P��K
 �0 �&�H<��|y#$^�@�%��1ޏ_2�u���2$%�͡[�y��X(��Щ����n����$��{�M�_�koA4wUI���N.���������(��hEg�bH�8�rT��b�i�!�JL��nF��r�������kG>�C�aQt�,Q�����2ۅC�l�?��- �:�՛!p_��婄�I"�@>T��5�w�����K���q�2�]���(���O�lG���^M"������h�ö���!͓ϳ��]}/-ic��Ȅ��!|,̛�6-�y��yk�eF��w
gƗMT5�bČ�B|[��V<�,�
w���;4&��n�F��?�o���-H���� �(F�l�컅Bizj���/���}��Y} [{P2�
�>� �KW]��?MM�ٽ�N���%�Ǌ{O���R0_,��gA�� rN�jޏ����x/p�������aZmj�u�EC���|�xCO㤩kb�>LU�C����(t���|�I��Ǳş]Sʠk��W�V�t�<RN9h3l�b��5�h(D��b���@4�pIam%�V�hk,�P����OF�4��LNxj}EDb��K�b1�.���yl�F%��I�a�}�0�G�cy	8���+�1'�(�2������ �L����Jv��i��0��i�_��	_�4��#��O�#;Nx<˪�ȟ�-{��*v�v�����+�G�V��P�0�3��՗S�J��Y��;t�����T�Σ�t���8�7�Z�[ �\1B�b��|y.
���}��S��H�����E1(�sM;l���m?'Md��E�A��0chP�^y/������o<l~xA�%0��Ŭ֤Ή^�S|h��<���m�*�C����*�{�Vd �
�N[7�-�
�Z$H������@T�^��c��[V��p�u9q����#[�z��`�]���R�TA�ֲ��͎��^��e���dk.�߀�JY��˩Fjt#Kcg�~�����2qp3�(��O��-'c��<�6F���v��?{�[��`I�k�M���֒<�R�щ�	��|áS���'�x����L
]��Z�+38������s���w�K�N<9�p}�7�����b��x5;�iqǆ ͷ�:��dz�T>�-s�:��Aܕ>6��w���~�+��< Et�'���k�������jV�΋�{3aǞ�%I��yp5��g�?��b����ʾP��*i=��3^�>�)w�����c&�� ��U��V#>Q7�)K�P-K�(py���Z���$JS��Ph�*K_�P���;�)1�e�`��D��#���н+[����N5k��z�����|ט��f(�u�?%���b7�
N�SN��U�
�lz�����g�����xS��\�ұ��	�Gj��<Pa3��SY�>
�3�@9���o��հ�/~�ދƂ#�)!Ȱ��w=�U��Q�o�탕��X��͡6���hH�����O\�0�)��c��3%���\m�{���R6qT4s���!Z�E��ds�UP�m�/�c�p��z�����-�)R	�e��M�Z�
�}�d��6	���o�c�ڴg�y��ձ��~��anPڏ�@��:��Mޖ��l"���xc�Yk��	�XN���~�W'��&T�Ew+����oлj��o���Z�|�L�2[����Hְ��FE�|�Y��'c��u��D�#cI��4C+ϱS��Ӯ����R�F|&�
d{�.��o"`�Fͪ�-ڡ�kjݸ~�+E�XuZj~�O�.�d��*��-�+(���/.W)��5�i۴���A�@���T��}��>�6^oa�,�; 4�g��ԑcA=O��c��,��VP*
4Q�\�"���W������T{ڿ�#xY1)f	�\X"n1�b^W�0]{�yPFڱ�J�ֲh_XA��Au�f�w���*�;$��}�;־�5_���͠C��[��WK��Ŷ;1aaj�!�C�;�6']zy�2��e݃�*����I˚�׈]+��֨���Q@J/�h�r��ޑ�D�-�C�/�FG�qQS�-.��n�8��K�� �S'�V��6Q$�< B�%~r�P���ݚ�ʘ��g��4��$���_����$����n"�#�26,*�7����U0U����DC��Њy��w�y����iI�.N�&�v�X�<������_/�?:�4[/�uQ��ER�6ϐ�"+.���C��cb���vY_)�s۳ �=�g@ �h=�� .�r�9�g��4�b���Jܙu#�l���^h$�F!z�]��	kd�}{�@��P���8yM��e8��_F� ���ѓ��ǰ\�|��e������j�7�KX��ņj^���:�O�#𬓐������~T��y�������}]��c��F�ma�o��3H�=�-����3��F�0�v�eߕ�j/�~�U�X5�>k�-=�n_u�V
5:�X$WI�(�9�U�x��Gd� t�샐f�yhC�&h^x�R��t֕PD@9��D���q�H� ��^��XBM�w ղ<#�}���?���!ZY�J��;m��k��L �x�#őͫ�޼":D��A��f���K�L6%��b��T�¹:τ� ��^5Ǿ��5���+n��d����
q��@��5SЏ^�|뜖������AA\4��fᜯ�?�Y.��꒘�}�(����e�T�k.�Ҁ��~�Y�(���}\sd�W��
��ע������_?{��>�`�߳��NJg_߳�s�tm&�����K	X )�2��hEqVQ�� (�wO���t��`�j&$�\���f��#'��B�uQر��(�)g���A16k�d%�@�^i��~��C��ܒr�~�r�_��4���a���90�H���<���8��V�m�c)��&��u��ET�4	vn���f�X=o4w#�oΆ�[�Qɓ׹U�����q%������Yev�����c�u1��`NM~�dE�-#���.�j0,|���5W�tUJq���^��O�%&�Ȗ�� �-`��駽 ���P?�ZTd���E�\�d�?vN]
�w�||�K_]X�&�|-iy%��¥%��OM�Z�Th��]���Yy���o�Vԩ��q6�$��!����hC9Z�y�Q��WܡG*&��мP^�a��ϳ�P�� ,"HlH��˼�J�(܆7�R�������f��?rr\Y���6�"�k�i�m��uޓ��6���)�x��ǅ�Ո5ʒF�yt#�$s��!hP��'0|����3zvޔ�vY���t,C&��}4�D2"�\R�N��Ɖ�9"�]��'���4<��B��_~��k^z�	��R��@�¦b�$E�f*)ʏ ��c�3Ǉ۶&�A&i�M��8�$V������9͞$h���ٟԬ�א��k��TE�E'����Ȏ-�L���c�Us�\sęF��������}�
-5|F�0�1��Q�i��>V>��6ݑl㮍�S��R�`�	���wA�{���0I��pG��m|>!9�Ui������3�/�2ov�+4�<�[��f����|�i���d�z���\�2�K�|�yY�n�y�%�<���X�!d���`C�YU*�Dq���z���p���Q����:w��M���_yf ~�,&��RM�#�D6^��f}�9h���[�V��z��U��-	9�G�&�:V�CKW���	z9�,��@
�{^�x*�]a$�J�0���S��~�cCx��^�dl�Y��T ס�������y��*R���ry��a����f�{�˵�Sn!|�[�;i�aA,��'Ktos�u̎YER�� MrgR���SU�1;f�g����7Y؊#6��p1�w���y�q��t��|�	�6}�aL�N�+>���/_�ȁ�
�#7&�U7�n+*���p�$5�TZ#O�m���Ů��9- �-C�z���"�&OgZ��&�d�%������wl�X�w�=3���)K����*��aC�ǙO!D3�T��<}_�<Đ:b���#W�O���[�D�L��[��2�V��t	�W�A�Q_�o*��T����B��j(A[EǞ"Qc/�	�H�h�͚U\.���0u��,��p�~v�hQ��H�N����)>��*��;H�Dhy�[:��^�ga�3n ��2����2'�Y��mz"td�!Α��W�Ծ�L_޸-<¹EӶ��}��`�,�E�M��U��O�%
�'�4$�۳�kN��2b��@�X5���-h�^�oԯ�ت1E�DI^˳����ySY��D��-�=�f~�Y�Oۣ���cX��K�Ͼ�,�SB{5c�����-�����y�v}�?�ӼUB�-��p���8'_�`b��Yr�{����Dj��y [�2
�WHN}�jØ����D�r�!꟫�k�y���b$(d�ȃ]
�^B�hp�dL��*{%m!9�[�f�:Cr�,�!3C}��>��D�SЮ5��L�%��ܸ�؉��	Fl΁�;��<������04�|F�Q�N{�Ĕ���p�&� ��C_�M�}t|��@�|,�,f^��I�^|Z�&�!5�P�H1-���Q��d����њo�j��:H�9��2ьS6�L�~ q�;��	u����x�v�/��E������`������ �y;u;s����� b�m�S}r$�c��}0�z=��g� �#Q�{$���G�"�GF#LP@W�s�e<,�� _� �"��] �����[�&�TPT����,�����г�9^��x���ο%�O�T|��Ң��x���n�v��҃�R�F���T��طX�.��I��@?��Z��zB��*�Gل��7i�c��C÷Q��x���_�x�Z>.����Nԋ�(=�Ǽˣ��;���*�堷���v�ò��W�X�B Y#|���ULw��ҷ�唒���Գ�Q�sy~�'N(�
��v3�C΁�O������2��	�G�&.����2_�A���SD���`e�2�L'�*.���X�p*�H/3�+�O�[��e��(�1�f��g��(����6���9�KO�Bv6?�O�i�T����C�lM��������otR:��AC�DfC�=P��~}Ro9IOB��������T(A�PP�о`0���xg�Q�ɵ٩�Vc�����]/�t�x���ߋ��'n�=�$����w�9�X	N�o���D�"{ߋS��ˏ�
��*�{���E3����^�]_p89�uv�r��z�5�Z 2�������	���ʒ�h+��Á-��!�:�>	��A��(R+*��F-����Gkw��� ����R�+S'[J�l��v����0�bFe�JĠE����i1&q�3�Oͻ��a~��LЙ,���IX�����=C����֢�`%Y��*�߭�=�w6g$&�@�?�[=�R�������z��o����0o�M0�P*�#<�{��:vg���i-R�V��L�rĦ�1AP7��.#������>vkF{�E���)8n���X������O�1-�������l4۪(1���'����o!�
���0�SG�#X}WQ���3���3�E���f�����*5���3
p�w���0 z�̔쟛�=����/�%1�1XO�a��o��jD���s����o�x+vCC�ҍo�.�}b��h7��TF<���kB'��A���Ww�3mr��Y��-x�OϱԄ��lq3���V��Q`�w��sdA��Ǖ��{���#�j6u�E���TO\����o��l;v��~�|X�_K���	ѧ�l߂>�Sp�����3�]�	�P��Ɂ
(�p�t�^s��T�D	/LE�\�8ݷ4+�k�������S�^���! 4���� �g^.�����x�z��W��7�����1���q��ʒ���Y�dR�?�AGr~�+���[˴��-ɷV���x
4 �ݱ��~ۂ����+N��	-4O��q�1��,?�T	q!��j�k0��Z���6��Uxd�Z��[��If��t�oz�0�<߉S����T�ߝ���↰�s����C�43��C|g�Q�0:�p>�z�)Y���𛍤�Б����.���Y'�s��y�絣\���Ν�j*�gdߣ��V�0a��Fvr����$�W��o���KH͔<�K�i������a��,��?�6~�����X+b��9zq��\�<�+�f6Y6���/�1e��]K�����-,Ӛ�6pK�(PZN%��˞���w��F�]D�e�6/Ӝ4�m7�3�
Dw;��w$��a����P0�����Lfe��_��C��W��
�?K�M2L�#S�!�I�1��
��q��I{��Z�;�
��q���� l�����>Gz ��MZ��pb
%��z��@��̆����Lo��羣=&���;��d����|m`A������W��b%�o_�Y�����?���
����][�����t?��{�~P�RF<����H�zB4��|��n�&