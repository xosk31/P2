XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��������_��qL�h}�
Ok�
�^�lEr�>
_
d�����TO mf9��k����F��y`&#�Y%R�͜��QC���3�h؍��Q�S��͐�7�$C�fp�݅ܕ�2���5af��`�&�z�G��L�jD���B�)�K�n�wD2��kĎ��H"t�w�ψHW�ٗ� �X�}*f���N}�Vc�>�x�c[HQ��
	�;��b���l����[�><@��U(����OJ�+F�-)˧.�7���Po�Z����푇e���Rb�קU�w�K d6�����yK8.}�35/,CH�k=��ځ3%7��ޙҩ;]I��\��7K��A���c| �6�@0��Vb����P?y6f[�I�u��M-�z2'�2k�\�II��{���w��N�|�*3v犈��h�Tg" �:��>3I���͑Նp?)ֺ�I@�K�+ K�ˢA;��V���ZИ�m�ݢ��<�r�[�{W�|���7�-�&
�Į/ٟ�Z@���ʪP?�E��;}C��}8�
K�0��4�����Ƹa���n�.1vp�fH�a�qDbq���BB�1�Q�v�n�)!d���n�X�@�Q}ٲ����6�����:{�c	����BUx�k�r�~�Y�ɔ�����^�΃�hd�[U�����^��"�*��)�&%-���#J�ǵ!]�����=H�7�cf��Sk;�W���"M�o}�*L�{��zmmd7O�T��l"n�l��RhWT�9XlxVHYEB    47d1     e90Y��izݼ�:�}��;5�p�� 6�ɽ���e
��#�I�:�P�o��T(,П�8���A޺��b��}Y[h��J�U��`�9���!�e3��jV'��ʛ��c4�]~�z��K;A��SC��a��~��u!��؉.�j>��:��gxI�I�eï��#E��pN���P`'��6�5G垮<(c�)�������z^_��(ꋳ���� R-�+�T�R�0K�㳠p7��ڜ^� �/{�Ԏ��/�6�)��aA:�8���	YE�6�����f��B�`��V*�K���>Dׂ1�\�r��0�h����:��D�@��2�?�:��iJAI�@�}i�̳�>DU���[+b@��ġ�w��g{�㍠uN,/����5��.���x���f\�+U��(��H���,
.��K���v��7���r#�3�DM9$m0�u�¶k����F2��ʈ��(��bR�{dp�q����^�n-��ͬ� Y�/ݖ���U@�G�O�Xߪ�Ӗ��.K�Sy�M�G��%;�lȹЋK��!/p�Ȏr#&��hsru6�4a+�-���/����Q��:�0xOᴜ1�,��%�,�LC�C�;�_�2��d������$�^�E�r��1����{� 2�`��ގ���L1�);�xg4���"�k#.0���<���B���j�ŋ��4���H�#f����F�3vy���T�wh��Aj�ᤱ���<Uua8mN',i2+��Ǿ=_C��T�If{������ja��]R��]$�)`G���A��)0_����ʵp`��| �j�����Wh??��:�ojiֽ����I0//����
)`Y0e>v�%�VHx�����k����SuJ�˛A����\�֡[����x$�Ů���8i	l�Dz�UD�|	�ek�m�@���RY��%q��f[hS��E��XU��D���N�!�e�SD)�v��ϰ
[��w�Q>�p��!q���tʸ� +��Â�"��:&��"U�"�*�-� Mt{�7����^wZw�
q�$��̋���{�g��:k����|�dyP�v�:�%K��	�;Fe�
�<DCD���i�}@�ʏ�Xt=%�Kw,«�1��?����O�4 |I�V��p�T�Q�c�X-�.��=Xȸ��K5CIB�cr�!��Kx|�.׫��J�@\I��1b���ײ�t�R�:�g�%�d�!���Ց!	V.V*��1�}�dr/��V��.��E���d��i4��XJF���������r�#
�$Gu�NT��/u�2Id>�g(��¼�1�2��K��|�
�nh�wxB�����"���H��s�jҶ'�["
i�pM���.�piP[�7=.��C��٫xR2SQ�.5"Y򑒿'��lje���$n�q��Otղ/jE+*�C��F�i���Є�	���`���*�&jp���$�;�W�s1:�_��6���0��B��E�jp�l�o�}��Swz΅o��@!�Ԩ=�|W�k	f���=ޫ���oN�"v'��852v�td��!�uZaV�ߕ�U"/��� (2W��;$�]W#�� ��=	��$t����LQ\x5���䴰�)��s1n�%sm���t�g��I���G��\^�71������'�q����ǽ��[�s���,(����E?[K�rky[�ʟ`���9!}���Q..)`D52��;>I9�ɉ��N)JG��v������U�U@�c�j��6!���ʘ$z+�b@�$A�`'��AF���`�s�UG"���GZ���vm�>�xV&Ka��A�����>���������$���쩟�ɫ�\�Р0ڛ7`���m_\YT�c9[�P�����8n?H.2\����w6�Q��:<4Z4c$�@m��̊��Ex5}ǥXoWȬ�,Fb��nt�P?V��BBr������b����}���1����L����f<Jv	s���_�܅�|-��ѐA�H*�b���U�\��� e��4>���U�Y��ĝd(��g�^ ��C�c�a�����.�v�t6+M����?4g�R$a������$/a�`Rڰ�A��^��C�ӵ���Wj��t^�+��Ë�L�B���#�g Q�Y\�uZԕ�T�����A�<����ȳsc���?���]~�8��!�aGǔ㍲�u�n�H�D���Q�p�~�h��$�P`�#En�q�=�ፘ���d_@-k�ˍ�;`���}t��)�qVl�xhOh��Ws����ҁ �dTT�H���Ҏ�c1.wiۖ�\ra�5�َ�ݮ��"z�My�h��i��bŪ bڪ ��V#��ږ9�7���R�NF�������E�Ե���s^�U|䤐M1��(����_Cs*��9��0�8�K���	��~(U-����*��A�i�8��GsB�����M��F (�-FF@G8�^�֮��s�i`[���B[�����|�~C�x�(��Թ��2�,	�1�\����J��0��i�s��J|n� �W��f3,��-����<�M��f��d2+����T�,�����I[p^����er2[�-��^���M"M��p��=wmp�U���g#�*��M	��)��"<��w���%}e+I�=c�����,?�f�U�@��d�q?%"^I�M�b��[A}{�9���2��^�j��̘�r�K4n��Ķ��撫��(�����]X������Jy�ӧ8tp^ �|�w=�	�:��}�`+,/J��	
�Ra�����OZ��<:�ӪQ6�_��8r��JA*���&���a����]��1&4cLx���Ӱ;�������\W��ޔ��*u#���}��X�!���2��U�.]/��݄h0h��E9yK`���m=`>��{.k�\�;vY�Q���*�u��ɦkO���%���kU|/����e{���l]������q4�E�/C�Lԯ��Yn����݅�.A+���n��O��~�6Y��u�|^�	g_�:��KC�f�Q��Fy� �����F��ԷVF�qe�Qy�~�>Ā��p��z'*�IF�h�.s5�<� ���F��{���/1���,D�llt�.�Y�d��_@�H:��W��)�M�*�� ��˒���������|PEx��W�-���(3�{��ң������d�{�9d��Z�����n��d�m��J9��r	r�_�u�|�&�6c��:8�w[�rS�� uXO���f��rv��E+�H7=�|b^�H��[T�b�Z�Ц%oX�k��H�;Ŭ���\�І���"3�e�c���A�XÙ4y-����}:nJ���Y�f�IK1�0Cy�m�Fm_=8��!WÙ�r'U��!P�#�+�t���L��-������g�ɑ��ŖA,1j�* �U\��pX��H�a)15���@F�O�9��)yӮ+�9�Tt���kb0�!Z7< $��LhD��ͫ�_u ���皕^Ū5��~�_�Y>���đMy���<�����i�'��`��o�e�����B�8��(x�Щr���d�1��4k�$i.u�*��z�Ck4q��'����dU49*��ʉ�f���� O���:KjӨ��]Y�=/�V