XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����mi( 6��Wж4�r*�ㄨ��|�*`�d�d-���	��k�́�#$ݣm�uwf�P���	6>H�Ӄ��Z���:ݬ���i�ԫ}Ft+�Y��c|�Zn���X��h3A��������]�V�Wde�ds� �?���L�>��5��D�ׁ����̓v'�(8��u�!dE���~�9�()��A�*_��K4~��ؾ��u��S?��џ� �8&7�ls��l1���$g$-�f.U����a_|�,wv	w�q�� ��iM!���a���jI��X'>q���|1GA���2���.PJ�L�i����L����d���.�N�ڕR�=�K����-�!�++���@�&#�]�/��;�Mj��<���D�'x�w#��4L�A��%b �$�"�&����Q�|#�u��R�~{�^���Ĥ4*ҧà� @��Q�ŵ�_��e� d�7���P�;���g��:Xy��lWƟWًP��������HJ�[B#�-��~3p��a炣��'���@Ǻ
�n�nmT�������0�?��]L.��Om����q�闩 �K!"�hf �r ��:���Ն6O�����r�aUD�v��A�-�pK7�W-�$ �2�P�-V\�e9p��M�[~�/~eal>�t���&C��AK>���Jw���岕�Ԓ�14~2�a&��1�ճ���߲.�딀�&�f�9Y��C�XC��T �6|[+gb���,�sS�?7%���XlxVHYEB    5dd9    12404'N��O������#E��d/v�i��Yf>��"�_��6�!$�>�d��;zS���ҲCh|(�%�ӸGҁ:��z\� �g��5P���b0̞<��.�^bY$����9h2�^��X�'&��;�$6$�T뚴6��4�,����Ă�׉W�:IBm����1�&d�C����{�U{̊u�(�n&��}�2h,g��/�pZ�1�IM$����_�� �|]��\>i�x��Ɖm�@� ���<�8���7FaX/�1TD���nM�d��NE�`T�@� �	�@��rI�4����x����еy����B��E�'V-e��HѦ<wTy�KفZ7��Ά^=�D4�~�'���5�St	����
혪��n5��/�%�
-�+	�]����f��*�.L��JO��VjjM |���9ƨBk�ߤ���xw�ي�Cĝ�V�; j�\�$u��6|Q==��e��zd��8���/�z�F��}-�|v�7R�1}�$����g77b��w���q�!i�S-�K����m5�ph�>�&����W�"%Z�Dpݗص;�.�'�.��a�Y�	cv&�N���.��C�o��rf'Y����D2�#�0�1y��\�S��[/��Nǖ��6��Bw�A-c���u*w�ش�_�2�9M��̟0�ĤݾX��a��I��R�U��_f�Q�,�/���?g8�mO	G@�h�jn�r��aҳ���#˔f��f�5�y�$I/w�3��B�6C��n���͊ɾ��B�`���{�θ�i��%](�CHs�����T�s�,b��1�/�^��
]�jl?*=%F5Ȍd�̴J�EВ�+��Gkڷ�+�H�uvI$E� �j'H�5���? y��*s����֝1H7MH�����rm���^X�1��N_�p��w
6����\���Y@�"ᶩ�����c������tG:�/����r�K�z�,�iB]�Pe鈽ڠ��fhehl���3���_���}���.;��B���}�np���)��۫\�j��]��7m�������8嫐P	R�@gk�l�����̂{p��JtGDX����jr��]�}��u�%���KyTfe 'O�& ��^
�C���O`Ѡ+�y(��U�N�r}!J�]�����c=?�vf1�FQ�]I';�p�Fo]6�mW��l3w�kO�{�5���N>Xm89��W����w7���h�=������*6a�W�t[�%��q,iuMo"v� ����7��U:�.,����<�MiI{KK��zK'�f%����ň�'���9�mVЉr�a�7�h4�rJ�z�� $'�:�qxӹ�F�~���H��r��4E�G����4t�g��냯��CšFA3ta^��E^��.��#֗�x��'��y������Z�V����a��D�9�"�,�s�}@�[�3
���Z��@V��R.��%�����>�1�	���,v�������=�`����daO���S/z�c{�[��h�^`HϢT��ŽEq9UE���o�a�YH��dn�"�B���Ş~l]�n�h6���x�q u�Vؐ;p���3P1]*I�Ct`t�Ѿ�,�48>��pH�x��l�B�vt�Uإ�\���s���������\g�b�%ϝÒd��gS�泣1���ނi~V	�g�	K,�5�7	��/�zˁ�uW��us���2Nc�W�q-��A�`��r��d�;9b$��A�$ꢩ�}���n/J�*�:�!��z:���x,�������ߏ2�؋��/��íŽ>�ϑ;����d���]�8�� ,ï�/bt}S]�{3B�rE��}�F��.P��4���uOwgFH�����C�YHu��0=�K�C��{��K͑�,�0,�Z::�8��
;h&��@��y�(O��]P�=7��y��1G�%�	Z�)���AA{�|!�LI��g�	;����$�<���Q481ʴ�^̐�K�$|?^gk�=qA6�r.�$�&��<�v%2\/�o���=��|kv��`Њi2̆:�q����78�n������Sw�4.�	]Zv�0�R��7I+�5'uZ����/9�gӞ�}'�s0�ᕳ�q���_1+b��g��ޫQ[D|�7���G��c<��Ej�cU�ﶰ3������Lh,��:)[�rZ�X8�F:3�ֶ"��NaWZW@ĝ�զV�W��lTC�L�b�B�<&R;Ǧ�\2���\]�S:��VK��_�?����]�D0m��2T�?<:�oЫ<��<0B$:&�� �ysRzf(l[$��5W|8 dZ�X.���Ċ9�$��B�.��^y-YR֓!iJ��U1�䘟w��`����	�e,�c��[%�_/&%W�	�ѣ�Y?._I�s��3< ��SdK��g��5���� �_:�`�=��
BU���>R#~-4Jj�##��������%C���v�ccX��ч�05�ٯ�/��s�=����M�C���°�ʖ�΍ICn|$dN�ϕ�ܩDH8�|8l���f,҅蚧�G�"Fe�w��N�"����6&~HbkfB~��I�ɭ��I�)$�!��e2���]J�:�P2���,n-k�L��)�M�䙲�]��	ס=U3����<� TK��ziz���X�`S�6��t�F�!T��F�N�M(�v�����Ёh�j�H�����:���D�W?���`9KPVӝ�S%3��]�б$���V�[ݝ�鈺=��3�i<� �B�����G��J� ���@����p�<�"n��>��D�f!{�25	;�$f� �{�O<T>���C��j�9��C&�X���
�_;���=9��9��NϤ�V���(�|��·��ڿ�e#�x'"/��@M�*�ظyB#*��޸���p����7�y�%�RGs��m�W��ع���~�V���(�m0U�읔i�/6�?Ӽ��9�I!u����ge�i�w�q@�G��K���Q�h-�! ,����~w'ӊ��\�Q�\WWT��M��a����W:��҈Ԫh���"��:��*�̈���^��y>���wˊ>͇Z�R�𷜋�87�x��<�R&+������o�\QG���^ܫ���~J$�,tDm�0�r��H��o��ca�y� "�-���9RG��N��ZX#cY�/�7F+y���������M���j�0F���&�y��OB��v�S�>6�r�:�z�_����AjڞT7��(�Hl���H�ѷFx
THI����M}K�R��F�h�ï^9L��c���A����ŬJ�!�'݁R7�vSR8��^CW=�ގ��G�=�ض�dx��
�m�{~�1�H	��}]+�L��ƣXo�f���7��^�rLt�H���L���i���񫙸}�V*��B�?>�ˀ�<��_�W�!�uz����g�b@�Y��@�2�l��xN=(���ֻ�����=!�_��Ć�+@;*L��䲇��������f^;mc�^�+�kЀl�s��"��a��h~LxR�$��T�}��y�CxO�S�k�Y�⠵]��Z�c'��P���(�i����qh���1�O�h�p����ilxÛ`��O����Y_�`�˷����W��t$=��^�6:��S]\x��L��>�`��=ʥ���-������$V��b���"W�Biɤ6x"�w�K��~M�Z�m��+��4��PݼgJÃ�9��9�t�u<Z�H�`��}{\��7��ĭ��RK���yD��Tr�~�"4�c�4{doX���+��9�O4���au���[�)7�7]��*v�^]�ŀ�>��sx�[t��&F�x!Y:B#�-�̈́�o�	�44;qIsZ��.Қ"y�/�V��l���Ԕ�|�@�\a�an�T���Elq�.���3O�Z،C��)fx����!�PVt�Փ��&�I}I��#T]HA_(���\�"s��a��Ϩ�}�����B�wah�z������nB��w�3�F����e�v��/��K<
���Is{b1쪩J+�Ĉ� Sn�s��8��?P,f2�ϣ�f>�-ٯ[~ȯ0���x�>����xз�C9+&�:���r��"�~�k��ܮgv`�fn)Զ0�um�pa��v�e��$�cC�]	H�q������������L�e)��U\`(���Lo��F��*y��jt����]��p%�5���%�2k��ئ���j�A�!�u�) J�������.�����͂wDcb�L7�9�����q�N��Ӄ6�|����҈J�z�0��Z2E�VMk讵"�"�+�տI�h�EPC�Ί�i�oI�Py��s���g�{�N߈�XB�tH���ٍ�2z�ܩU2Q������ǈ��2��7&}P�5*��\�Aau��l��� r�yJ�y���Ӳ�?�=g_B�@�0|7>@����E��`��,��A��C(��!��/��+��S_��\�zf�\�L�"���{��ҫ�k]��Ϥ)6�*%ρ�&Y2�����q�Ah��> ҈�E?�7�W�|%n��Ӵi��:˩][��Dt/iO���i�a�1_��P�R�&�ZW�9��F ��m