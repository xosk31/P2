XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���)�����X������r��hTz�U{*	�<�9���e�}'H�,�/�^{=�#ԏ
�c�% �v�F��Q�_�:_�3�i���K��+<� E� ,��,ȋ��_<����HΓIʱ�������jJm/��)��
�5tƷ>�$��R����'�j�U<�\��./�!��iD�O��(B�C��_��$�q���Yu�d,zM	Lz�#a�v��?F�i�u�T�8<U,�[8�x�c� )��������5 ��py�-�wT�t���G��>ZX�h�i�1
B��G����U�wj</C�H�#��堣hB��۶~
�~�^���dT��6ߨ+T����Z�������1��q�d�Ê\-ç������hh׀e�@/�%'E8KW�U�傶�5/G��o��`��=)�>j��a��m���:~�hXa���D��Z�,��Ə�8�Y	"Zk�� 4���e�w8����Ve��Ձ�bMٕNʞ�u!�ⅿ��hgo��Ŵ$I=d�¦p�l����]���k�%My��uJ�������	��`�,�!�����Kv����MSt���O�<Yrw)��$jm膒����g�1����_�wBj?}r�a�zN.Z.�ݧ�*�b�q��5ɳ*op�
'$3���F�N�.%s�ǿ}�>e�m�����,��Z$�svAqn�%��@����N	�����湎�F?��[��}׊�0`c��ι��T��2��GWUJ�7���ѬY+o�$;�AXlxVHYEB    2a4d     c10���2%��as��+�҅R�HK��H�8�壙��r*sp~��9��M�,k ��p��F'[�@'r�Vd�S�o
>x6J	m)uU�u� ]1(��_+<�ZEk�Z��q�[I��!D� p�&��:K`�������&`���M:ys�8�X�w,��<���V�䚔�҃���H��k��n/
ʩ�h���I6׹x�;Dԇݍf߲7n'E�����Q����\��-6f���!�����/�\�-�7�M�	�W̔�@�>|˳�-@Z���r=w	tG�����)d��j����60�?Q� �'�{%�T�G?Gר$|�����(�ExwY��HK��	�Y�+)17���DNA���2P�H�y�+���H���T]8�С@/�E����;�7ls�I!�7�5���59:�4�*��-�׫�#�{�ȼM� U�$�M.���>8��7h �P���T����r��J�KߺNM��;��kL�ٮ�*:}I6h^4 ����iʩ��w|�]�I�+�	R|�& �ܑ�hS��3t92��^x{�Aq|�U�T�E{;�Y�G�:��	t�)P��i�{���],k*(�ٳG��bT}U�q@�a��mR3c�%==~�i���ܩ�*��o�}0m�:r o=kg!s�0��WM�fȚ1~�ݎ��WrV�pF�d��z�k���H��?��W�|�{�rxŦ������ ����M:�
��t�̌k�cxH�K�?�7�Je�B�i����RF��R�6��~�VXT�\�w�����&eD�ot�e�Ԃ��r�]��`��ŲF[�g��Dj]��?�2�꼐ze;�|��n)q�agO=︂̂#D�M7�P���7�l�_�Q$e����o<l��<u��z����si�cHHR���)͸o[�<q��L>���W�ͲB�l��S
U	��k�uc�mus��
��;< @E��2z>y�Υ���6:�~fm�H��.����W��#�#�ъ2�m{���	���:��5��uJ@��a���B��6�R�AϪOvN���2B��$:����d,����K�A�"��7�v�``
Q�g�Ʈ�)�������$+~+`U�f��	AI��U9��p�I"E���j�=���s�A�:t�S¦�l�����y�7j�$y��4fƹ�kz��읭x)Y�G)��O�]PM��Ff���p8 ��x���a���Az�� z�ix=p^i1�%-��4�~�!������ .D?��)}���g*=��x�0�QC�$��m�9��(d���[�����>DB�� /p�?7��LجT��~w��+|IJ�Is��E�#D�K�7�$����D4��jHF�V=S+����T/i?�.��e�iڼE���,�I�V��'�8=���g�8K��F�YQ��M㉹�w��h�xX��6]�Y�8n0_nV׈�a<��eO[��U��i�K���U���0�����Ʈw#]�r!`../���[�<Ljq����'�'��l}��'>�ćM3��s�Y􃱁�7�{��~Y�"�@@�.���:^�ew|��~x��P�N����իQt��'�.n�h���H��<��!���F�]�ň�]�8��[6�����*ŕ`��qСO�/V�`<UhF􃮡6Ձ8N��^%��\�a��W��T�� 㐈
h�Z�R�U�p�/�X��JO 199�Af� q�~�ia�~�(R!��oe%'����&'��a)��E<�^;%(_D�w	rHx�����$��4FQ�a$�%���崿&���E�5�e��|ɤ��q�r�wSO{�N<}N��8}��A��H2�$"^mjg�Z�}���x׬]Z��[����@�h^�T2;�Ǌ�I�7Za�$9�����Df���^�W/�P�if�->R6u����ۀK���F���qe����x��rIK�>m�<�!d� f�|�Wb
�Ɣ����8ٲNʀ���9�A���S%'L������Q��sq�<'aIbPoS~�ze#�مoz�sM]R��q����!w[B�����K��t����&Z�a�&����D��)pq:�=Egч��Ƭ�֭D�G�����Kn�IWA�+����U��˸7��!�Hc%L*����TN����0�%�k�+�D�;�x3f��T��v�Y��@3Y�!/v JGk�l�(��Q�?�9��@nj ��#羹sÎP�s���϶�l�s�ɍy))�p7�N�]��0� ����$�M�ԓ�����'�A���U�v���9�@�0	k��]�oF{�(�̿�y8=1�B�n�.�L.����n�QA;��.Eg)�d?�Z���a>o����������בk���YT����L&���㣪�~,�5�}��:�h�a(5y`i� ��S�^Ù���-�!�W�~��8���A�7�t�+U؊�{������F���^��W�$�B6_� 64$�W�U��K�����u�r��vu߶jBU��/I!��,մ�I���Ԩ�祸���&˵m���+A���&�E:���|��`��_�C��Ӆp/������3����"rcZ�y��Â������E��܏6sz^�Ɖv�R�L��:a�b #f^y�]�J�s���^� ܇�9V�Y͚-���u��%�߫��ȭ�:'/d튽�3����"������4����}p):��E"����O+S*cM{�����H)�R#�s1�U���+Ů������5��\3��(��E�;q�Wi���j��A\%���`r�0!&w!y�h���7*X�+��d�b�����΍΄\1���~^ح.řM=��5C�^�ds�n������V�h�h�c�\n�Y􀈧�8p�Er�?��|Z#C��NC���8�e�Ң�RG����MI�����U���S�:������t��7s�Uu���UK��jH|b�^���N�Q�q��[/Y�g�N��� _t��Ee��[�n �@����3�	aXSP!��䮛X�Z�