XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��m!�tm;���&|n��!NU~MGJ�gY�4M^nW�O�7~S����q��\/6��7r��<U�^�!�ރRYў�����#��9�W$�V�n�.΢F���vwq7�p��s@i��1����Ql�g�=w��$鳒��Y��Jf�3l����P�U<nLG�,�p�1Z2�:k&n���zF�7݉�������	E����ȳY	/��j��y_(L�
%יݐ�/�߃C�`ww�Ҳ���s��8�6��"�m�l|�=�mL���^������}0�W�B22��Um;��҉[�,��&�)�3��ii��k8���,i6	�H%?D��ˆ�xS�@�A9��={�F���<m�u�u&�T���Ǿ>�� CƓH$r���R��]^2����h��q7a�U��e���$�o�U����ۚ�L�iP@��h��_�T6=?�]4���(���sE*�-?"��@dn�3��M*��`�"�Ԁ�<���(�ً�Q'1�"y������L�B����T�걗��� �ֺ�L����%�~������̿x��L��0/ynF�� ,�߼hI��7)~xG���*.8�X��58?/�ަ' �1;=���7\���iS�%gxvb�p�g�R��t�l����&~Xt8zKf���I��>�js�l�Dm�'�v��)�	ڃ�����9�����"Y��t2��X�m?7/u������!ӷ럂�=�V��Hy?�`�Am���ܶ�J!�����=�z��H�<* ���XlxVHYEB    fa00    1f70ڈ`�#Ҵy�/��-<�����J�5F�F�(:��İ�`~�X�Um�jo��F��-g8�t�M���oBqnV���v�(� X���;�&�������US�S	Ct���D�����k6��WvS/��o�@+�:�ElY�"5�$K�/Ф�'�X3�P0Kx�����[�9�Tg\w�)Dk�c�҂l�x��y�_���N����l��A���a�A�m��-�?k�������ƂRj��\�u�B�a�i+>v�l)�,�:�e�o
�����[�6΢��KQM��|������5�Y���4������t��\b[ٛd�p�Ư�ѕv2���u.&]i;h3�X��G54�WWQW�+�,A��T��`�tЪ�[��1z^R��xY�j�e5`���������q⅁2)����a� �h0�@�n9�~��4��Ȕ���}Z �u��G��(���U��(G����tH��8�k��p3�E�V��� �֨�V7�/#9���Dξ����[B~'���l��9ވ�k$�~�!ް�ۨ�`�U�@�:��V_�3�5ir�Ěk��6/@s�FOB	[�'2k'3x\��mO�p��[&���i����8�OZ�^��'ٕ�����fU�G���N��$G�֭���7*�vw�����"-�������3޶�;l�"�G�� ��j��$�c�Qt�OA�Op�ȗ��� �f�ūn�Pex�VԔF�9�'����Q�
d����&���ϒB��� "')xS�� >5g[����ݛ���۸%�蘧�'��	1�@�)��Į���Bj�q+��Lk��7��44y��f=�F�Q<����Cm��u��
�{&=�<��s��0V�9�c1'ʦ��?U']�Q�и�a�6�Nm�oi���kb��^�DxA��^	&�%8+�xD�� |t���'�5��Ɍ!�>�6�Ա	�������J�ƿ�co�PF�xv4���= �	LCFu��g��#�)���G'eS|�$�L�$����
}n���V,T"?���C=E��"��͡a��H�x~`<M�Yޘ;�hq�� �T=m��m�L2�SؽV�𾏗y[�������s,v����J�2=��y�cV����8k�b%��yw?�%��)��²X'�ӉZ٥�����á��OaW4a��:A�ji���S��όt������w�o'�Œ�$�1�.�hVPN%�XǻՂ���P0Z���X�I�S�d�)��h<d��'�俳Fa��^Yp�u�s�� � ��8>֩�[�p���T@-!J�:�c��tT�A	s��n�1�x��P�X�c�lY��W�s�BJ.���6��+���yx֩u��Q��<wa��윝A�~,5��m�e�~��H�˽���Cm���������G8�E���=��W�0��geFb�d2-�N�������1R&��D�/����Ɛ�����5e���Z� �o2Q�@�|D��o=�"��E���6^�����Lb )4���:�����*k-�EǸ�N<�+kJ ���)p?Ggw|/6��Bm<뉭�N�κ~�-�zƔ�YH�%O����$A����vA1g�ns��{$��
���h'x�]���!��_��J,������;������h'�i�97����y�&^=˲8�챠W�<S�H${�~�@|�UT̕�F�3q�d�TOJ�*��xy o-����ل��M�#B�գ�W5iZ:�'��?wh���u��bi���#GIfV\���I�����4�Ԋ�r?^��叇=��p��$
��w��y��
�U��˨ώy�0N����"�c�r�?�����x�	Yo5�+�;68��x�&���;���Az�x��3D�V��x����$yv�l������\�����b����<�P�+:��!/�+����9F�ARN�j�B;�_w���V2���(��ӕ�6��#<� .�����Ŭ�2Cj�r2��{NT� �u�m�����2B0�a1�D�J�R���U=pE�-7��������
�?�d{=7Zأ���Ӆwϑ�j��H���0�������޶��^(Uµ���׿߲�\p.W!Ԫ�mV���nG��J�r�Vц�+��sV��+�d��	札�Ҹ�J_
��>n���M4��n�v�3Y%���<X�����]ε/|d5i��"��i=K
b;@�*���ȵ
���#�߇jo�G ���I��;A���;�̥ʪcǞ��� �>��t��TJ��ų��e�}����0�*��B����Ϝ{#.	��'"5x���6p��XM�������}��P_:0�0b��#��%M�&��A��� �|�F�w���������=�,h���T�A�v(�A0�ч@SO���$��Q~慒���X�)Ji���g�}l@�
/��W)	��^����?��iv�,���'�T�0��/����~g]��:� X������&5p��gJ�(��u�o6��Qm{���C ��rVIk��	�Jo��������η������x����T��L-��V9[]BQ�Rz�[i}uK�7�tQ�������J��%+���"�H(¤r���˄�:X1�t�G�F�`J������\�_y=]l�6T��� ���rTe����d�f>M�c��Y�H���\�NǓ�Y���uD֩��0^R'VT�Sp&D
�jy��q�C��U��+�a��Spkʹ��$[���IO��~u⦴��R�
E�O�ܓx����:�đ��7�X���?B�Jh *$FM`�ְ�����H��g��n��vZ��$��.�wцV��
��x_���Q����b%\Ö)�c��;d���8�_1��e��es�o��a�� s��F�c��(X��؀��~	�wiDH��?q6顐Q@�]�>�:�u�v=��$�>wr\_.�Ac6s��%�y��`��/�h�Q�N����\�r[֫p�mN��ɰ-	t�0E�-�u��!bX�ˊƊ�i���źH�L,!Y�v�D=.�"g@����K��,�=[<#; �8���ʬ�q�R�4��So����I�B��S�8��>�A|@KH2z��Za�C�
�B�r�?qc�s�Z�g�L(��5�%cse����d�?l d���y%ɩ�UԢ&�w��I�X;Bz*: ƚR�f�SG���s�/��߀�<���ְ�ךa��F4ꖲ|��3���F���s��d*9C�0 ���V��L�B�}��¾��r>�����Unx���@܂+y�G�{33W�� ~"����t8�y5�'�� Ǉ�sl@n{Lj$qw�q0x��0��A�?���*���>�:�X�
�$������oz É�톭�&��
G�,r����&5��ƒ[�`��e�IH+����i�K*�>J�Br(���wT��xg�}d}o��{`l��Kx$b���̭��uE&w`PoH�F&ʽ��5��5-h$�6�1w�Кr�N��5��S^,��~X߷;�Ψ�W����55��M`���M�����I�e��{�v;8������ n^S���v�$�+u-�]�����C�eo	-с�Cg0q ��{����]�:���Wα�ϐ�~}�,0�n|�A�M��Ii�Р���~u�f'
B��S��fėS�J,�Vo�@���O�*�JgXݥZo{�����04ϸ7�͝�^��>\m�B�
���ɠ]ﶩn�O�PX�P"��q�>��lv�V	��q�W+a�쏰�%00Kk��K>J�����j��}eS_���7q�Nڍ�S����)�ܻ��c#�vt���9��4&2�f<z�`�i��B�P| g� I��vU�zz��Q���t򁏕L�0�Ap��u�s:7�A��hO3����FYV%[Q�����|U�AOT�U��1��/mcB(��EV����6'B��˜�{H��V/1[Ty���)�t�d��*'�n*�6�^�/����G���H.��6U�e~�f�!���>jP��p�J(����H�6��b:D�
?�}�R�7_jO�5� 2�)���V�L�'E��mU.1�#�Ӣ��&�}!Z���2��rKN!�f�t�|}k�F��y���Z���SUz�A�W}R��P����3nvp��V���q|�n����;%���z�8���z�L�@����Q%{e%T��3�eS��vꞫp�b�����x�ɻo�Ӓ��Pc�w��^���5��M���ͥc��\T�SFX����!
���)��T�}ZŃ�;#�d��+�'���Xʇ3*��q)ݥ�E����]�f(Ba�Hk�J�F38)�,<~�c�RJ�N&�P�z��A@�^�cF���_n  ۖ*��	�0�5HFrp��&$��Wr�q	X����z����Ϯ�l��w�����Q��>����a-���o�r�z1��cB�������N5 Q���b�O9�`�����˒r�~d�P5ì�H1�㣊��6�<���Z P�hZ�> ��k20�y��!8oԤ�D!k���KcǎoP��y����[s�҉6k��4�Uz�7����g�B���1u�>����/(���'ou�6����1��x�Q��ޙ:�GL�7�%�g��leB�!��*�4������_�Eۿ�xDQmgVZĥaބ�L�����'����B� �12a�%c���~j+7	�x_�pc�`�~|�
���YYo��O��惩ϸ+�-�`�1%����y�Pa���ߠ�T"��Gϴ�eo@����=ޠ��v¦L��a-��t�E����T�id
|�Q������Kf A��zƋ,�l?8�&8%%������I�ᾖ}:
����(�X�z.�:��J�KUx�eG�ܭ)C���q'Q��bs6SZWVo�^{���Ah�q!��%�k�ݢ�B7�E3�_���+J��M�W܉yیJ�g���Y���-4����,�����涧��5�]As�&C�������V3�x�E�hd�O�nd
Q�T���XRdA2,k��������(��64^�UM�9?�b���Ơ<$�;"Y�w*F	Ƽū�^����^sO������I�:�����E����L��x�c�,�J9��������G@*���Vh'��s����PU?�F<[�o���Ӕ`;��n�5n���7,��Do�[E�%ױ�!e�eEQ�\U y�fk��4 ��8q5�v�<2g���:cl3R�Ij��Ys�xVu�p>q���{M��|c�zܔ"�� �s��4R�;~A�CP�I�F����cL��oe��J�A#E�>��!k��O��+3܂���%���9}��"�eI�U��W�e
΅��e�x���\ci�XM1,�M�c��r���b4���W�20���`6ZI�L޾�o����lr�c�R�l�]�w]��F�#c���2|�oD��{��D༗�eA
$���c��.����{뢘�5���L��|X0�>^�����
UH3j��o܁�)P��ԌYX����7:5����|1���,��$H?�ɌKvY29IM܁� !+�d�Kn0k��Z�]�f%�2�f�ذ,]�gL]}i<�7 i�|�TV;+�1V��mAY+��T�5�2S2S7g �
ԉ9�"�c�ܒ�+��0f�~n��4ɺ�b)�9SCq	�4�{�5�$�Dˁi'8� �k<�Y{���_�M@����\����3	o!Ip���N�RF��@�8���C:0��!��v�wktsM�ZF�<Տ@Dwg^N��i�i�����\�[U�ů�v>_I����Ы%��BI�K�����(��4���a��3��{�@�`���}I�L�I�yQQ�`y-�׀��u�k���\�]ђ\H���o�*�ڔ�P��B��^9"�����v�ro�I��j�ȫ��0\�v�r��Ift+/trBׂ��3cX'����i�n�v�5Aۚ��y�֏m/�[mԛ�,�M��,�c�_lޥ�&䖆�	�xh8b�V�3���琫�z������|��h�h25:XT�UU��Tw��/)���J[ ��55��H�}���L5��akK�����ݔ�C6.
n�T�#pO/�*%��O��ֿ�t��+Xa�M��i�&�{)|\������ϻ9�L-!S@��g�J7��N�������.���vK��0����Ş#|?��2�گ�J��6�}K1�m��xC8!k|�h%����Ph� -�:0|'8Ki�-�2_Ƿ=I�{�	e��}q��<�6�١���pl5��v ��.y޾�cR00�&.��8�%<�� ����u�r��R�KW�s�;���jBH�ov�^w�:�Y�t{�Vtt��h�Gb�-��6�'�Ke/6���cx���u����y���;6Y(A���EB�ϰ(�-��^��pV��FNp�f��*u�j
ahG�������/m�"���"��)bG1OG���7��V|g�L,��䱹EP�Kx1IR\��������TJch�?��5����7�D�K�(�a���TȾ�e�f�"8�ި�=hf��\ײԼK��;�̎)D|���$�#��	�2�_i��q��x����	U{0U���:�'���Gʴz�._4�YR����!�zu�� s�<TQ�by�6��M�&�e"�zp K�.�9]*��z=��rȸR��l
N=��Z%�zmץ|�E4�sGΐ6{6�Y��8�bO��{H��I��b������{�E�DBbK�����'��F��ģ?�0V��������>&m�������*�\@]SW轶蝮#�����M�D�����t���;�<���p'T�-@�h���D��͂���L��Vk�?�&�f5k�k� }�!	i�=<�e����e����w������R��������q�T�]ê�-޵�Q1��z�-�@?�$�s���C�l��cH�W�4[ν�T���Y���kh*C���m�����
��S�{g��'��a�A;XbK5�T�6�]�V�=x�6��6�6�n4B@$ � �؛B�6u5h�ݣҒ��T�ɅÌ+^Z$ٜ�b��yD*n��}ʤ�AIf�F`�T�/���W��v��2��df6[x��?��mfE�޴Dq��f'�2��A�<�q����
ф��U�����0�J���&�Z!�̥_�T#yv���+�؋�ư����~?W��S�5���_� ���`�nZ\4[9l��ƿ��zG�k�X%��LP_���q�?]w�e�x�{������S �w�5�ix��~��7�g�i�����g��v����OF��D��z�m:�<��?e7��7�=���" M²��?!��3BZ���5���i����iG��c�(�ˆS'���8d�V�In�/�㴠��DF�Vl�R�v��.�a����p[]�&\Z��vi��7*���٧x�]�K�P@]Y�c�X�8(���+
(��3	�Ic$��3�gq�Q射�h��Q},y�A5������ŕ>��GT�
�\&��D79��c���sѸHN���F�9xd�;pK��i���BTpI����V����
�r�DMm~Wk�ح���PV�"�ٔ��.`�V�K#��8G����1�-k���d��\O���.D�����_4b�w�ށ�Ǥ��F�j���fe�J�6�oIw�f�G/>��81�6`����Z)�����v�k ��ZӁ7Z�N��V�� X�0F�����" �G�����E��@�:�,2kb�+|���z������.��:˼�ʞ��r�����d�Sn0ߵ2��v�>���:�N$6�o�;�iD�{)��+(�gW��"�C����ʟ�,�N���d��,��ߟ�XlxVHYEB    fa00    10c0�G4��� ��ۭ_�V'�7k�hZ�dy���J�����1(��*�u��52�m����Vb,��ld�U�*>{m�u��s�PK\j�.Y!�'�l��2�y�t�J��"~;!�o�O��b�P}���f&ڂ���g	��ؙ���B�.6u��hi�B������fXC��oK������������Ѳ+�w;�����������F�Vtsp�')��L�9���%�м���E�m����_�Z��5[4�1f�ʙݗd���2�yP��� s�#��� ��<l�w������Gd@x����.u����D�1J��[�	�,("�c�t�~� `ʊI]��F�x#��*{�<��j�1V���A���6�;�a�����x��sã��,{?z��M�9YG�dD�z�P���?����\=f��>����&��	)O�\� 7[w�{H�� ^�n�o�=] ��'����mX(O�t���Bj��e�9��M�hAP����zũi�
n�@{f�9�{X9��kZ�ˣ�?3�i�rZ��>��fz�H�a�@���ĺ��ޱWp����2#/�!�O��^�6c����O��~���S�]�h�|'�bf�d��L�t<���w+��j��y!���;�C<�aH��P� ��C�
�b�7s�|<Rm0����u����.��%)2�h�Gu�&z�!�n���pvW?#��+�T/�p0���dX�w+�8%�$�������9�5�`�Z�b�^�)gZ5��tr�S�=F�j>�JD�6=pH't	Žc�<�����4u�8�L�_^FڂE~�[P]o���?�1�^%�cs�e�=]ۉ��UO`�o*=)*=� � x��ҫ�00��d�L_���AF�A��XV�u�����Hqj���h�#���;h&����&���	]D	LA��nS���Q�4B��T)V�����=�/?��sG�&�UȿL����|�S<ueK���yI,�ZnA~Dm���
	��FS��G�����m��^zM�v	����n��-S7p7�س|F��@�=7�)b��38>g]AT
�P��T�b*���7P�D�tr�$i|�|����lAg��	���8�B^�-7,[Zp�?p��kj�в����6R9����4��_n����
LHy�@��"�i`�U��0��ʤY�3�!<��,K;:
m^�+ؼw�1:
�eD�Hd�gݕ���	%�#0�s|CT���;��cS��2tt�����(>|I!��͒�zW��5�%���7�2�N����ر��%s��O��r�V38��9@tG�Բ�|��e���y)k0|*��Ԗ�`���=��0v��ٔ��j���ᇇ�k������K˝-
w�:���O�]*����$�\6���C��0�Q�����fEP��n.؋2�� C�E� ^�������p+\W�]��C�k�.K:g+\�¬�����Dք����\����nT��6��6����ף��~9vWp��+ęhs�z�u
"��C;3v�� h/�K�h���}�&�\	d� �az׺ċ�7Rm�25��?2�5��&��!r.6;Ո��)d��n�e%ނ&#?x��7ȀM\���p����`uN���@��+�3;B=����D����<Y �#@�5BK�hs3�jnd|g��hVӪ�Z������Lȩy�$0~��w|�R�M�F��u�D�9�.(wߚ��-��/�>+���@'� �C�y9�8Gp*���R���
�?R:�uZ���*�Z�E88N�T8��{kC�],"��L�Ff.)5�O�}PmH�1���sp�!޴�(�&r���.�������a�֨Y��sw�<��5��^�Q�$�(�+G�)'}�K��#��x��3��_���,n�*)b�3���_J��ඌ ��0׆��G�,-s�a������a�^�i��#�O�$c�����L��yPcQ�`pj����m�[B�X�LR��5&������GXм�)"�t�*Ğ��6�ai����k"8$b�>��䬺'�P]�T9��=:z@T�z�W1_�Öo����C��u1�������T� ��4����>����I��ϘS�5�2��W������ �8��F�?��>�8�4��m�zfWN�x�m<��UIX�����B\.Hlz/����b�]+�Qus�L�ʕ�<{�~�;k�8���N����B���^�Ն��?ЗAY,�^�:-_�Plm�(��&N�7��o��.��`��B(�Ύ�X8L�jS�]�I9�9&c��/�a^�u+�h~^�b:�r�P�=�^�r�l��r�sF���۟���'��	���j�ҼK��P�ˬAd[�V<�Yn�?s>If�\��6@X���.3Wf�V-6?��e���"���P�Q��Cņ�R��$���؝z�.=��.��p8<����^?��fD���d��u����sS��x��g�eha�Op�]�:kk��5��A���ؽ��a?7$�န!�7#ǐ]�w��z8:f�,��<
�g��R����s��1:��z����T��`��,��S5��������SB��#|����y9�>�8�-(R^M��I.�����V���<���2>�ib�7�(wz���W*tR�d�V�cBK!C��E�I\3���I.��$�x"f�rZz�
��-��ZbK�z�ǷÜ��zY�.{h8���5Ӌ���K��hn�&D��3�����Օn�`����a��d3T{���)|�5���1��3o�)l�9q2I�}P�oi+5:$[jY�Uɣ	�PF°RK�˙��YO����G�8#q��T�!�㇀.���Q�����>�ɗ�LD� 蕪�9�%��?�l���܋b�L�^i�fQLo^ӵd���Ib#8;5v��]��B��}ܞ�:�l
�e��<�ɒ)~�?�����I��Q�>�1#���Ű!���I�J;*��C��mYW�|>a���N��-3��F�'�Y�w�-}8�3Om$�S���лM^�%��q�CV��LwQ��&�+l���V�9���X�}G�JJ��`��!�<~1p��7���ͧ�SI |��v�`�/w�GĠ��"��C�#9��O��|?AiM���Z k6QS[���h�e'��L2_�HZY+�c�#i�s�U� �pt ��:+ңUѳ�w��/�?�������j3m(#��0ϩ�e���`tt�`)���؈#qR�^��/%�^[��@�(rz�t�B,\qi��㜁��P�ܙH��<���aLn%�Ѩd`|}��{i��a�
�N������[d�YH����F�yA�h��ߨ9�s��*���CaU�b�fQr�v� ���z_nB-�dd���(�rȊ���J���A�,���3�a8�˦W�O��b��89!Yv�2frc�G?�v6��0ɾ�	��GkKz��Bt՜�{V#�6�Td)���;��A���^c���z���[[��mV��T������S���1���������3kE��a��Q����I�;�<z�0fGt�o�6�ـ�dY���;�ǏT���WT������ɍ�{�t�>޽h�(�˫�i��s'2����_�Y��k�@/�r����/�8`��N}X}���+OA��[z2�q��^��jU���TJi�N��}Q`�5���(���JUč&�P�6�n�_�CЄ��V�Z����Jֹ4ڢ�;�_�� �V�f�֣�� ݭ��N%P�a�G��#c� ������H��C1�;���Z�U�|]�� U�w�"�J:�щ�{��c�W��q�'HyAv��ncEb�K�
���e34T�k�&�@Y\Ti:�H��ȯX���|˾ �,w+���3����`@z���0=�����&�ln��fʣ���v�?e֥}����o��n�c}�D��cDa�tVL������t�?Kz���l�B�'g`�I�]Lz�G�|g�(���G������P%�e@2M�;��s\��O���N�ysIP����iaiƁ��g��{����Yf��pE�Yct͘"�"�����e���/T{؀�=�g��w:+d�ɿ�1�;�2HS���o, EcNed	��1�5y^�Ѳ����-
�ߔa�ab�A�I9j�����5e� iϗ���Et�S+ҩX��O�����R�o]%KWC>�����.pay�(8���p[��[<Ym�XlxVHYEB    fa00    1140ɜ��]���ԫ��Oq�.x��3���H��k�����yQ�UG�\�L�L#$Lߠ;ʜ��EI섐�L����D�(d�)��W���r�-�S�u~�U/�!�Y��ٔ�o��k��Yj��I��	���|��.�y��#�Kw]������%Ѹ;r��.x��SA7�\�0�W�F��<x����^�'_�
-oUJy�x����"Ӹt��bcQR%>Z&��2v��:�w;�1W=��q/s=}�/^��E�+u�Nb=�&��-��?�BZOI�}�B\'QlW�w��c� �
sA�Y�]��l���k�sQ{�vhԂ��l��A�:h��e�y�5��"uz4
Sw@ՠ�BFL>��]���K"D�-;��Kw1�nDN0��9�o��d���`4=)�BeT���Z�fyEi���J��!c��Z�y�:[�Up����&/�p�_����e^~Y��\B�#0`����9@L�;[i�L�0��︧���c�x�GH�;�p��ͅ�F1*�Q.����iv���.����	7|�`�&�'�x#�������2�f�gd�z�&��	��˨L�/pO�ǟ{�k�<����)�����3�F�~�rgg3!�&4SO���!�J����/��ѕG'w��ܶ"�`5l)Px�-�.:�J�>����]s��h��*].��a�=է�9l�%�s������dɌԔH}~;�*'��/eq�J�5�P���kv_��4 l_6�6�����i���<�H��2���� 
�,�C�6��Ł����u�$�4��E%X��T���*2���^��0^C���$Sl���T|���Կ�E��Q3�y?���P��j��:Hw;�=Fg�j� <C�3���`MU@7/Pv*��s��'xګ��b�2����7tE���6�ӝ�\Ɣ�M[�*���	8�����"�='��ĦS^5$�~k�*rG�+KE�]�5�N��]�򌒕���t_\��AB���6ihί����G}�ٓ�t#�����h����8�>���%әNb�1Dv��r@�j�	sE�}~���Hϡ��.e�i����A%
$ĺ��|�`U�(z�).FN��U�����԰�K@��_y;zR�����c�ɢPL��`�*: z?I	�����~I�3����^��uC�L|Y�o@�jl@�ﱳcaԔo�zw9�X��g�c]�q+���%���f�dy��.bD��}œս���5���h;�����H���b�EB�;�m�-M��5��5a�%7��3[�N��e�.?�8 �*U�ǜ�F��a&s�#���T !w�[7�Rq��ƺ��ɮ�����@B}/���+��s�	�PD�V��� i{�<��2,@����SD"�����E͐[� }��a�.�ğڵ�ݼ~�!�լ*�� =�_-��,���*g�M.�lVa�����*e�GY���?\G�y�݆�FcX��n���"7�!�(v��:E��!-��av�T5l�����eT\]�6?���{��D�'�/@@��vc��crʅ��y��)��G�k��l�����5�z�v��!K �\5���,�KR`5�U��� o�v}�u�n�}����<1R���n�m��i��j����3 ���
�܃��3�o�1���e�,��6��Ѿ��Q�2A.���$ɐ3�0��c��*$�6�E.��|�%��B��B�4Jj��9� &�oS��y��'���n����e�Q���=%�i�q���mFZ:����e�W�y\lL���"�n�C��']v%��y@Ëi-�5�2����V8~p�������5Xp�A_��&~�
���S�~��-�0���v�Y�U&6���#}�l�B��8y �7��R<�{�ǟ��'��_�))zS��-�x9��1���cg�H�nOb=��;�e!�jì}�PA��RC��|��)*�f��8Ƒ��m-T�Cb]K�����tX��)#܁�!7"�_he���^��M}��;eA�oNd]-��-��v;N��:��%1M޿��2E�\��ˊ+�s���Gr����S�b���#�U�B�4�݌7�:�X�DrbT\@
�^��W�[GF������e�#Z3����J�kg�p	/����|����x�~���K۝�����.|�t���Tׂ�J�����߱5�1�n�߮Jk<��
��*�*��Z3�1��Đ��s�L&i��s����x���A�L�A����#M!��,���%W7�q�597�#n����N��o��p��u�	B|F�x�YkP8��P�cb�֑`A��S�I�=��F[i�E��6���$8�C�Mj���j���k^�����Qc��x60�@F�QO����]���<@$g�|�B��w���5��{�����gҕ���X�OM*\
���m���,���T�����/)2>��3�j����C�8a�u�H�X��6*���C
!�d��6�BvK8�br\:ulz#�G�E_�kp:�kL}ڊ8��X��Y��5���K���r2~�h�7� :�s(3껛�(���L-�.�:妨��*8ː�Z���,�^ת��_��cK�K���ܚ�N�o�_V�d �N[+*���q��'��	��5����ʙ�B���ZXj�s9�'�\3��k��-��H��}N>�oS��5�j�(����h8�@
�F��{� ��dPY��
%�ҝ�W�}&yh:��5=��U$Q���I���{��M��P��&�N�:{9:�{�1؍bq�� �ςI`1�����G9Ip>D>�3������y�k�/z`��V����2����<ą�(,�*����p Ҟƶ� ���կv�T��l�6d�SjkZӳ&ǿN��p(ШR�~~pT,nzQ���J��3,2�ܷ�eL�E���9��L��t5��`e�nû�� 7F@*f0>�G3���M����5��o�5.��[:���=iZ��^���S���jf
)>�gD��}����ë��35}'Mq���c�ܵ�U�r�"�3�,�Xe�S�e��l�,�U���I�����:���
	b��=���j�uȱK��b�ktO r_�|������$0޷ O�b�.�I�b�4M���ۉ�X*���/���I6d:7D�a�b��~�VN����{�S������}�����X<^(��< P"��JX��W�d}8�������k��������΅��zeÖ��� h��դ	��J"9�`_l ������WtTI�z�H
��d���G�b�U�q����h+�<*�jF�f�ύ��k7p�۬�`І��a8�w}<��&�ki��W����>�7��Z,Ig��A�j+V<�ko��8��<�z��1~	�g}K���d��O��e��:�hI�rI�xa�hK��!$�	0���~�zo̫�]j.l�%�������z��.�[X�x_$|��K~��5�h� �9�;���^͋d/�R����y|��O~�k�ی�u�.�j��� ]G�
Ʊ�������*��x':��ܦ+��ТL�<���Tp?����Z�ơ��]���9�{�{I�,���~|�9���[ ьf\^z66��L,I�Y�J��-g��=金#��N��	ISL!J�e��
^v� 
�I�}���e�{������gL�a.VV!�3��o3�鈓r�wD�KȘTǠ.+d�^	�%�o=�A��j��0mHm���?�|�t�W��z������P�l~&ӌ��H�U�����B�B�q(��.X��>7+��q�3�s����f��+���(5N�n��c�fq�I�	���&�!���S!Q/�˨6KeD��-N�q۽<'Y��\b�����h��m��P��[=��ֵF���g���^��+M��w�4�*�c�H%�H���bn�#az��;�c�
�
c��P�3�𔕼\����cN$�/}�t�yu�<��g �n>���+P	���)]��߲ʦ|��0�������U�'�X��.�{���U��D�k�����n͖?�Hp��*���nb�r=+��Tv�3.Rٴ+��p����d+���<2�E�x=$P)&|Xe߭c�Ӫ�.�K �\v_F����6+Te$�>ҷC���|��!9ó����أ#�:�&?o�r��:d+_��h����l��vci�����w�ii偝��A�	��'���IϾ" _�՘1r_�`p�	�,��G��<�0����
�>�(yc`"?�0���ٶC��3���	�3�و7ꄏ�^�$����~�B}�n���p�D�`[r�ZD�cRl�W�[XlxVHYEB    fa00    12e07��:.��|�yƧ|Z੎��Cȝt�i��ʀB�L���?A7H�X����΅�v*�[G�!k�V��L[��;9�Z���R M=�_�G@+:u�m"��x��1�����`��$2�*Nl��ڐj�Lk�H�R�v��>0gƛ�(���u0��M����v����;>�,qڃ�P-M��B ��ٶ1�V6���EX�����ǿ.;������B�9\w�+������h��2~\�s]�"�V4ޒ�l�x��e�էԎ�v{\�Z��\������䃘s�T$��zێ�&Ƣr+��LO�i�Z��NJOK;d��op��Jкډ��9%�8⽻����DG�z��J2ȉ�]Z������{)cފp�zR4�IՃC-D"��#�Ap��=G&X�U�&S�e:���T��?���zB�E*"�?�"�� �H@�b�V'��]��?s�n��6Rr,���Yw{������	�Ԫ��a�a'�^�P�!�&�53q�u��$m �`b?�(������x���>��J�*��)�-P|��,h挮3��uhӒ�}/+�f��{�a\ޏ���}���;Z���B|'kRC
G���|-�bص���G�uH1��L���[�a��]{��io����L�a3g4�g|$6/�\8.�`5���Ȩ�����-Ĝ%n�'�b@�e\�tl�_4�� �C%�NMkHtYpj��'�64�&��Z���T�D�k�z�T+��[� O��<�ʲ���kj�)��2�B�i�y�`�#(%andŃa��I��~e���3\�)��#:�Q�n��m��^:���H磳d�uCy�R���d�}s���t�a�h��;>c���-1ƚO!D�Y�ko;�4U��
*�em5$���F��y��XNARPT;ܷ�1�	v3]b/�7W����[��V~�9p�G��\2�eY��ʂm�V��GM�O�Xk��2vȣB�z���;8%��Ki[ nڠ:��CT��n�QI���L;t�3��!��E���w�4�er��؉F~,�n����-�`�Ӱ��A������ԟiY�?����_��gG��S�j����}��)�(�{���8�ޱ��Ѧ·8s߳0�������:��&�����"i�l�u�Z�3LǓ�`F���������Y���R��^fJ	�W��E~A@2�������j����4��3� �f��u)�Y��M���d��o���R��O��|R�}�]�ɶ����S��ӕM�Y#��{GG�۔���Ύ�PS��7G�q�Ǳ�ޙ���*��˴I�tɲaQS��/;/�[��S�T��0�1RMh޸��dO�Ϥ�� ��~�Cӟ��� �Ĵ�(�����<⤾;�7�ܽ����#YzHPypY~@��n��j�N�F�u��J�D���&�fn�*���T��IF��g{���'��kh%��k���}�bC��N�3"�b{�������j�bl��̓����y۞�l��K�`ݗW�0���k��S-�;E�"*s/����z�9M]��G�ϝ��l�_�J�VlM���_�}闿pw�ZNs�^�x?�/]�o�9�ĳ@��'ڞ)l�����@�-��M�n6����x@�/�N{�����Xm�X]D���h��(E%�:�"���n�#H�~R�!w�
L����}�������"���a���3�4QK"���G���T8ڄaOj7ꃇ�;�OW}C�9��K��E+�Ή9:P-\��ǋ�m_M��++���'ǌ�c��KA]Һ�%�@��4;�u7��U=������~��r�`�{_�Ӓ����ZhjG�/ ��v
:��pTrD�-��R٨m]F)���U��o6i낈�zf`�Y��p�O{���­���?t)����B��%��'.j�jy�QjO~����D=� �N*�N�D�ؤ�xo�N������~r��Ȩ��t嵊t�)��.)/>1a�c�M^������!B�����/F������3<��H'�jC����m��vM0�(:e��ĭ�JG5L���2�-B+7h4����Z��������i��m�#�F�7mΣ��R��C�گ��g �]���Y��)�ۃo��+�g���f��WJUV���[0ؐ7��@��婪��0�ԎQ�˭,�[ā;��Y*1������!�"H32;s�L
L���02� ȍ:w�I�_3�R�O�/�i���,X��*茥*�U������ͱrJI�����o�{��|7� ).��/~�3WW�#D"�%ݲ�u���r�O�Tp��q��������x�/L��,88�6_��@w��7*H6�2Pc��r�憉��%��K�ò<� ��(b��:��<́D�aR�@Ij¯Qz�`9��a�CvR��kh0�9hP�Q�.��g��l�MR��V���@���E�� wՊ������-��&IУS����D�R��7�q���e�
Ss�%�Ͱ̚u���uSuJ�n�:/��F79'�A�ά*���*�}eTF<��Jqᆩ��B�Y��oja��{	�#���ɉ��d�R��6my��i�����YҶw���c�ͷK!�pnU��t�(��edt�y_qص� ����C���nȋT������#;��2α6_�_��=k>�TZQ��;���[%�n���	�29���1�ݜ��26M�KiXZ̫a�<���=�8��S�yZͰ�>ڣ�E�h�L��4;��O�)�=�5���\��v�0�#xk�t�M��<�jAUS���S�;��O�- �Y4+�U�.����`�|x}���+O Z���.�V��һHi���\퇕R7��S:��y_�������py�ɑ�E�8���w�CWإ� b��47Oh����H�iW��N��Ã8<r�K� f��~��Br�󯭛p}�[|���U�+O���k)���V!SA,�L;�;��K�Hk�ϊ�U"�˛˴�-c�L=����^�Xn�*�2H�j�9��v�C뷦��[��o�u�T׾eQC��!L���9���� 6���)bB�hހ?<j��yK���_��(#7q��D�j��`����`�[^��)��!*��*�w&T\���\��-�E�vOw�&��z�q>��X�o��bG�f�K_�c���G�r���:4d5aDhod���s�ի�"@#�)��rʏ$���=kJ�C��z�p��]�0��p2;Ik�%�5�iæwO1̂����v�I��i/57���j?�D����W��a�F;��6>�����ie�����!?�>�����m��ЛivXU�rl�*���U'�O*�Uڄ�S� �@|�y�SU�d�ɸ�cO���_?����}��Ը�[s:�2uEO���އ6�-32k�@v���K;�꛲ሲ�Q-mx&J��ݍ�O��zkLr�o#�w?	�瘽O��[}�])���7�y���7r�ER~}�5�F�R�����C9��X�4H끟�{�\1�l�!i�b:�BP1Z���M��+�9u����E\�Sn�0RVfֳ,2�����f?_󊐔�}2y�Iz����{H�o��.H�j��x�P�ï?�$�<k�D�:���!�y[ջ�
��R:�V�� ��খ��yz���FI`�����]���j�Nqm��$���M�ڠL�,�JWY���Ǯ���ʬ��AHz �h���a.��c�ӄ�+���@��������]�O[��Zg��k��®8b���{���d]�W���ʜ��#XU@|ߵ�H�g�:T�K�Eq���d]3��)WT3 ��`]�Sc��6�%''%;k�\��[��*��0��������/٪��h�����Rż��c�9UH�U�y-�V�Q�� %e� �з K�C��d�I@������!*�@A3[��I�PUDJ��+�T�OT8L�`��OI0蠁��8�4_�g�P�΋������$�*QB_}�ȌΞ5t�P��0�v�N���ŠK<ȇ�d_��5���	�����@���x����fdl�@�Ψ��6N�6Z�pg1��]҃�����R�\F:kT��bAdn���܄�i���ھ'�"}a���ˏ�@�z?1��5k���잫��+6*��CU�v���E��|)��f�=R��O�������<��H�?�v{)��BF�z�L�9$E�M����z�Lȁ�=9���-g�,T�6�:-O�`���h���3�]#n�!  ���q�ė�7Z8�����)ˊ1�R��f�A���Y�k�	}��%ԈC��8��.b�bo� �8�Ђ��>�2�>��um����8(ː�o����Ma?�M�QzV�������>�g� "e'D�.�q��e:[s�\� �"�^��Ԟ��b�)9r;]��5�����P��`����px5�4�%���z�ݤ�p-��\ s��wU�#(�A��P��O �]��n��8�#�2��R�A�`��ӓ
��M��j�6e~����-�W�sS|@!n�0�0��ׂ]�1[��E���(	�-�ĕ�s7�ά%W�U��,�0��L(X�I	0��S�A| &���.����}�Ā��؊�U��;���[��L0._{*�����e�rpEOC$�f���(��.^��:� ��r�qI�[�o4�*�_����8�d��f#�_�;�"t���X�d��ę��I�B��f8�CWT7�Q
,&D�֯y�(���T�V6|�d#���>�*�Sx�ӧ�j�����GXlxVHYEB    fa00     f50�PJ���<6��i~u��4�P��!�4���s����f�$	u���g	�U�p�w�yk�4�d���܅���뽭D�v�)Aµ�ˬ�f'�N��:�u���Wu�g}���/�]��n�hF�W��x�-��2j(
x��X~!�gR���jjF��Ul��z��+�d4�Y��W";�s���sU}��#6ݺ^���rB�N�hf&����7�"s	+��}v�5�l�>�gk�s��i��y�GN�t�!��9��9�,���f�E!c ��Y�q請�>L ����Jq0�邙ɉ-���6��/�.z�\��n	L�M6e-و���(Gsv�)�f/�Ӌ�q�y�~�������fⱥ���.�.L\�8���$f��o��n��x��~����C��P�]ަ@��!�@��V���Ay0�·�'�wY�����/h����)�$V�[�~z�}$M���$�,�-ލ�$*�{����\���Ԁ�&Uf?���FA��*��Db����ߺ��A�Vo�����8������6�!
��<��,�,K��}*ѩ8~��V���9�Pt�nw�����a@���Č��ܫ�Z��G+e�ڔ �
enOJ�����g;�N�T���Yk�H�4~�h��6�w�Z:JF�`�Z$��US��!�"â��SŬ�e�)XWP�0w6!N��&�A�r�����6�I���tO��ɭ0޴Y����*V�-An<&R��б��`v>�kJq0�|��r���'{'Q	u��K�(؉���Zp�?�-������,�6�r�Vڤ�?����`ywA!Zlt�b1�n�đ��WQ,�uD�o6�m���Vz��9eb j���9��v��J$(���$}�_�O�s1���^��U������X��&i�% ���Ody�*�^%g�=�5�����'
�74�+vj���'���S���|[�A����G��6�2��<2�8�+���N7������b�q8s���ihUm�j��Ȟ�t1l�&۽��\!��iaZ��u��S6r�0�}�VOV ��ĉ.�l R�K{���Dָ��?�r�(���&�s8�LȘ�{冼��Z��93�Ь0��[;F�ܨ��wR���\����wE����\H����j(�Zsb�nZ&���})�n��$��a5[�}�8[Y$túg�=���5�xK����Ş�h�FIx�W��g*rp|Z��J�F3�"�E�v���'u�9��iF'�+�:�4�G��-�k���;ft���)�w�S�5ZXa�U�ы�c��`�����R'�(��r�H��y�8�	���$s6��|d�W�;ְ�O*/::f7���gͮ6iȦ���g��4�5�X�Zx�����:)i��芮��S�}�>~��$��[�#yۮރ��iW�)�C��x�RX5��y�S34�>=1c�=2���*)�64�L�bA�?��y���T~�p�EF�W#��Ԁ�]��7���kB��	�0�#���;�/�(Q����#t?�����޹�I���So6��	����b&�sQ�u�K��n��d�F�f�6��/|��t6��q|1�5��D�zď��ܷ>������b3�S6Oxb��Tڦ0�+��A��咁R�����3f85Y�e]F���ٟax)�*2�Z�!G�����;Z�;W�R�CA��:&q
�3�봍݊.|��x����rM��8�H���`�mX��X���dB!�@F�P���3�*P��6n���8�F��`Κ���5������G�e����ԇ.��i^ Y��N��у����k2h]�x���m��anb�!~%2�kM���_[+&��>�BQ�A'����%z�u%�B�a��:�,ZG������,�KEHn��ޙ~g��T��$�U���:�-����rЯ*o%���j����ma����Ğ��Đ��k�ͬ�t�Gؕ*&+����)U@`C;������5�q �r��,�^��]����Z��Dk%�^�hLj�>4*�8'��=�>�|�:B��Jd!���1�ؼ�N�n��#���u�P\G���Qx� �'=g���y�����׽�^��
��2��3Y�ݔ�ǂ���%�`u���ߓU�lp�7�{�*v��|^$��{���	⠺h�w���IW.���e�_��;|�}��{�ȞIR��&F5��\���ݥC�&q��	G`s[�&?�����0v��jgd��;�5]�dS�ch�*�0h>(�4sZh��t5@�6�w����C�����a�"o����O��=��#�OsF�L���oH�i����wo�NF�����m�P �8n"L������x*_��1�"l���B*�x<d�?����X��Z���y �ˉ x׀(/q�S�a�^�������q���k?�%&]cߓ��"H��hc�V��W��
^�ud�Po�'D8`������9t��%#<�����K��.00�\�5�ڼ%�i0��.�P���<}y���f�-�9�u��Ԝ� .����M�k��Tؙ���q_K����,�ٔ���[���~)�Fɶh	B8e�|
��s���U��P�<maм��.�0Di�nl����@�=����|i�dD4�n�UU�Ƅ:=�u�.�|�jz\��m`)����#�v����������P�#�*������i����a��:��O$q��gn.�p��vs(U *=N("���p)���L9iw�b�]j�Ɣ�,�&B�I���K�с��b_x⍷��9+�=)U��t��ÂR�n�-�)�l(f��R��{�w�������
��~�0�[F�[��O�S~�i$�]��?D����5=	q0T�:�%lMQ�M��6�����R�S�S�e]�cC���"�T1t0
��������Ia����iG����	%8�*$����	�R�5pb�`�u%��LQ.;8U�>��3B=����*�M���BQ+���N��][�i�*p�l�q�#f6���EN�ݟ\װFf�0�;�P9��k�^�S�w}9�r?�ꔫ4�v�-��	tQ�%��t�n�
�t�x����_�	�scC��z�����!���O���B6&X"k�[�#U�GA�����N��1��K�����Y���v�N�(.o\T����lǆ�9L�,�:]٦Z��|��R�!n���XI0E��ŵ�4|��� �B���t^R���[���$&�8sm�5�}J�?���í��Bh��u�!���mb	���p��Y�}qdԩ�S������OnX�`F��'^�O]�=�I��r�+Nq�2�"t)	�燻�^=cN���6'�HI���jaLV̻N��)������D���6��X�AZ�k�R(�_���`8�QP��M+��w���)O��68��Tz�Y��B|���o�H)ud���5���Ro�9|�f�0��V=�S���9r����X�o���֐~����f˚��/�	�4�p9ک�%S����Q)��9%�����r��-i�!���^��D>�66����w7�D${���j?�b2k��M����K�f����q�#[ۃ5��~M�Y��'}�L��b�Q��h���5��Ƞ�u�zs�(ى�y�9;�S;¸O,u}{�dߢ��ܴӁ~���</X�^V(]|iJ�6`�
���+�Sr%��V_kf}����K|�ބ���ox�b)��Q�;֜�Q�h�bJ�r��]�t�3���ѮA���`_ʴ,�ר��"ٳ��Y��/�S6��]��U`�[�	�/.T�g!�#,��$m�������5CҚ�|���|������F5&���P?7��XlxVHYEB    7273     560猗eB���<���.��	C���������;4цTV/�	m���ŋ2�:@+:2����#�N�xb�b
��~��	���=��D�[�"-���NY�bm�NG+>��k
&�bA���0�e���Q�/v1��� �c�9��mFG,�w<��5���%6�N��6r��5uYQ���ٜ�R���ܻ�����
�]�es*on�����u�5�קO^�G�t��bH(}h
'ay	����[ڔ�-��q����{� O���%��6]�8Ҟ����d# f���Rɲ���Q /�ىD�W�{�=i�	|;ǐ�i����=ڧT��3Rt�:0��ӻ>5#���m��jc���S+��$�>���b�R�d�P$�r�w���;�CK�f�9�IJ�-:���b�I$>2��RMt����&l����� �Io:���㭆�8v��iEw�^&�Q�-��(�)F^�ݵ��������fC(m�?.nV�;��F�ҵ��3!�nM�Pњ8$�������W��0��-�
��!�K��J6�W2c�n#U�I�/�|#��[�
�b&(�L���,�0X���+O�!oNDU,c��ۈ֯����/<{Q{�!J��C�����5e��J���g>R��S��q�1����_�NG ��A�X�!۱n'�UI,,�'�h���l��f��/P�dd�$�A`���#�H���|������ �k�H����_53����4�7�|�C�jy���
ɿ��	���h���r��`��}1���j%���RY�0�@�|���PN��s�i��T�_�70Ooȵ|�__����w����!�&At�dJ��#�+�\��b�[�q�V�K���Y9B9���.��S�*@�Q-%�GwY�0�J5�V�\����,�t�"��k҆�1�G,`Bd���7z���B�1��.� ��s��+������D��
�*��$����8@�Q�co�ދ_�U`e�U��;�o��b��O-��q%E%�"�w���`y�sb�]��=�VU��+b���=-�| |�����R�[�\�Yy��F�8�����2ȗ�Y��D`f��c�g�����2�GWr�],�!�h�l(�Is�Ƭ9��c�� �Ο�����|���]!�\L�X�:v�ZՒ��ӱ	G�����5i� Q�&�t��~�@��$[R5QD�'�P~N5E{и
K|��Cp��Cje�*�m��ϯؕӇ�ج.��[6KgQ'9>�P�0������P�i?tz5�~�%j��A��<�컚ߕݱ	b�/�)%e���@�� X����rD��W�j���q`�-�t�#�y�e9�i��h�Y-�