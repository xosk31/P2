XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��2�ˏ'NI_<%1PE8�a�`Af��o�yf#~��kt}BFd����LU ��c��.ZP��o}Ks�C�П�*��vxgi��2�Z�m,�;��� ��Y0�֡gY/�~�ei�Ѵ�b'��:��u�[����R��
�3I�@�#�KP��<e7�1����Q\���� ���m���͵H\g}����[�W��B���ά�6z�a(���6����q�z[!Ar���$�}��N���{�g����)�T۬�32RI.���~IVv/�4#��0��m��Ӽ|�w�E�����<�}On39��q�'^�"}���>�/��1�6�%��������W����f�7�''k�9zх}���Q����i%i�}�3L��X�0���k��ke+������^���(��ʧ��M��2R6��c�\� u@_7��ί�̧BY�?񧴆Әʼr]f�*�S!&�~�j���+v�%
E� �2�����9���&a�_�|�o]�Ru���c+�{:��	4���F�,K88F�vo�q�ŏ��n��y�xk�B�}�N���soS����;Y����6h������)��D7�z�ΐ��	��E̷æ��Q��[tK��W�k?9*�{��n,sN��
�*����]���4Ş���_V-��
;E4�g���c�r�H�݌b�؂���T]M�˕#���ځWaps��S�Y�ג���}^ch�%u'�ϫS�&�=;-)ܫ#�e~�m�̴	�~Yq
���^�l$�`�XlxVHYEB    66ed    1670�:=��EФ�5g��<�;v+������E%aQ*�L�,��o--|-+���?�M!u茖d���'Y@K=�ZwYP��g�d��>3mU�NHУ2�r���8��h��54=�F�G^r�{�����h�/D�c���:���i��
���f��˯�:�G�>N����≘����}�,��'B���?%����a����y�,X~\��=�X����w<_����TIb/I:�;���v��D=�ē����kA����Q��%�C����^��
�Ц,���޽J"U�(�B`Z�%N��3͂��Y��-���;��L����_����ߤ��u6���&�@$���u�x8���9��
���J�S ����(!�2#�,si�@p��;��%�˒�ٯ��qݴ;/����y{��p�'�ЏnF5�G"�K�H����)��f�Q��N����\��.��.y�wt������!E|D�����Ct���A� ]*.�,�k=�=���~g`����D1�f�w���d��lw�[�K���p������ז��>���U�ܾ��H2����Gu�mW��8g��Y�Bء����@�#1D���y������Ro�,>�����PR
����x�(Du�`��hv�.ۦ��
�x=�.t;�-U�,u׌-p��1���m����tN�`��~�j�V3_ls~�8�䌷z+��-J�*���\��#�o���
_G0�ƆD��}#8�R���L���LQ�U�4r|�O��ş�O�j0~+Zm�\-����,��1�=���Ӳ�$����<��矞���O���?s�>�%��y'P*��YK��ĉ�9�rV��m&�Q��8)�Y����(D@׾J�$>nx�(�J~Ī�����%���x�X��H���1϶Ct� )�_�uz�D���U`@Auܺ�����c<_y������&���A� �n��ԭG��)c}�?��'G����"#c�ШO�#��Xx6��.�Ά�fȤ��!e�gx�B�],��]0������	3{	"�I�Yx�P�����Gԫʗ��s��I���E����a��`dLCN���vO�w���b�Z�VLQ���9�k���u����m�.����=
YP��d�M���-�(��i�/�q���\z��� V�$�l"���	F�g�2t���Ţ�C�����:�z���y ������S|Vɻg9� ���w���^�1��6�Gd�#"��.�R�v}H�tx�[��pT�l�JzoW-h �+�ؽ�>)(�k�e�u[��\L�K�.�;�Y���Ux��_u�{Ӭrb���m0�|�#����'H�9'���;�Zq7��'������4��_X�~�7�������I���Э�C5��Q��Dt�qf��B
��_����wݥ��������H����i[�O����B�UE2��)�>�j�71'�#���mJ>�2�$¤����o���x�h3[g��O�������"��+�OM��L7�q�u�m �O��l�AQ~!�s��zdj���>;8B=�'����t��ƽ�;��8����[P�I����9�{�|��Oie#ԏZ��o���Й�ǃ�X�?bB=*F{@�p�}ю���T*|w(�f��ň���U���O7v��A����a�=�����Lf��*&8?�m�+���,��-;i2���ٻ��+�R��^��X?�W�:!-��Vmw,?�:�LX�l���y��|`�w��?����ʤ6�Q<--z��Bwq��������J�E�Y��륃e�$F:��)q��n�J¦�yj$��%~�"dlC�/��u���&xQ�� �5�A��77��g���c遠��
�ޚ�eX����H�����Ԅr{��H.����2�l���8J�Cria϶�<}����$�y�@8���͔N�u{��糧T{��������#�7S*��[��4��z�z�\���^�GQNI��t�4�e��x
#&�e;� _X��\f�����@�p�~���u˨&`��f����#�0�u��>R	��vOz��"�3�[�և&ʳ�7�O��(a�P����@�d�؉�\,���UW	s\�'�����4r�kxB���������F�����a|�U�@��{Z����`�#Z�60��Z��'d����z�������˸*�l�O�֥�iW�:�ei�.����ր!�8��J<.!�`�v��`���z9�,���|�`b��~ێ��e�ڷ�bl�3�L�1t��e�'~���*~��,�,De$�O�5#��v"P��V��@$H����k�ze|ӛ���~�	 ecH�H�0�a�bB[�K�
a��������O]xsGXxmɧԂ@�!��x�/�!lQ<��&,a���o98��xfMKs��a�D�7�iQg �T�@�V��ң��g�IVCw�śPTq��]��т��[_N��,�}���ޝņR˯��<!�N������$���
�\]���ybo-�8��9[��J���6R8��v=��B��?`9���*���$\,1����4ń���~O��*p�, ������WT*���b��A[JEm�$7�MƠu����rz�o^�!L9j���e��+��{�kڣJ�@�浽��A6f�?��|Ȩ��Q9�p����E�ʳ cU�;ޚ��Q�9�~l!�nʡ���Yn���WɚX�r=	��a'm3��/�"�7���I��6�AwD.�����4�n�$��x(����ɗ�S�H�����A>z�c���Utd���w���a�5�u��!+WI^'��̐����Z��Yr|\=m5<)f.�AO���`T�.��X�2�����لݪO��p�r�c5
���}U�Y��d a7��"m�7�T�m�|yw"����\E$�7쬃��%'��ZAe��$;�I5��R�Eᛡ:3�[��fF�& �i!�$����=��A��wԘ?w�u�xh?Vs;���V�����&���|HZ$���B@��"��4�Qqo�:g��n���H
���<N�փ]/��D���A�s$����:�ˤp���qy��4�� �]3E/h�y�3� ��U���28*]�g�a����:�#9_e��&�K`����'���\7F�<��܍<����|�+���l�!-/�Nx�?m*�Yt�쀲�n��(����c�?>���V4��"#/���7.¶<�.(��vcq�-2�g��`�����6�$��Y���5l�!{k`�`�؟p�zĉY�bu���]ΧP�	�q� e�G ��L��Ț����nNcZ>}�۵w�OԦ;�`�����3a�-)a�M���K��[̐�������<U+�
׳��%/���PTK$M� ���A��
�fb|����}�ֵ�q�,�^�j�=<�6�6��^�m	��|���1U��$_/��h��;3&!���ᕎ�>���GF�n��Å�M�Cn@k��X �c��ɐ�ȴ�1���1>�G�(�A�D���1cP�Q�#̒E��d��J�A�8Q�Mf|��KV1�Ԯ�}4��,3<�}5�]9�y�Q/5��j�;IfgpX�Kw�PǢhkA���A(<���s~s��\��@O���V�F'�_�ߴ�С�~��������k�n���@�-Σ2G��WK�U����[2�HIb�?�ō�[&y�wz�A�I��(-x�@���&S�<�'��m�w/jA�C�		~j��N῕ںYh�8���� )D�i�z�U����C	/*:��c�[��7[B���`Z��4b-
1n����,�꺡�G�g��V
�Edq����4�d��g�I����MR��J�j�f�� W��,q�V�yK�qܗ��Q�3;�7�3��^i3D�{2s	���)0����5Z/A[�j>��������8 �T+����d�6mPh��`.3z������-�Yw��ю������oj�~77�Wر�H��y��~��P���>��9����/�0�X;H%K혽�a��Ɏ�N��}��XA�w�#��ſPu#���F�ŧ�)��go%Rt�+�R�C��3�#�(���v�Î��.A�h��'o��[Ft vy�4�	�.�Uq,!bD�m�(:RT$u�a�f���)��2��xZ��2e��]��E�g".1�w�ds�MFH���el�h�sB�r��J[(��u�?S4j��ﵩ���� �_E�e���d��j�҇"�'�[6{<.�ɯ�{w�II�&8���ھ��X��� �Ë���{t���e��m�><Q �N0D"�w��q3��M>Գ6���!s����Pl�G���S8��=z�i����CJ2�&����v��!�Qz9R:܇��!Go��3����5cdhO�.�A�E����C2��j�s���z�&��(�)���%4,�p��Ti_�nv�<�8�	\��sH^���B�E���
G�?2��Ө-X��VLw�>���oZ%~��/J��a+�*"At*.*|rv���6?�mn�z��ڵ�x�#�J�f��Rb���K�S��n�[�O�\�>F��a��^�,��J��e �`ՙ�=<?B��$g�;kC-y���V���ںLuq�m����j�R1��B�m�����c�j�|Ӛ��	����=WQ�+�b������I�>5�02q+?ҹ��M��`LE~���U�5%Euy+�5�����c�?�&lS��N�rm~H'B��z��`����0��_t�KZZ��x���[���@m0[�� V(N���0��C�Vp[�h��;Ce6���<"�e4NC���d�%~I�r��<���w~mx^�Q9x~�C�+F]�=� �.yD�ڲͰ�<M� �R��a�d�"�G���� fWն���_�*�"y�W� ��. Ҁ��s�W�u�w���}CgtO��J�M��B��C.�G�uT�B��s[xo873��a���-�����s��!�gR�đ�5;yA��)E3}ޝ�t��Р�}��Ѐ��H�x]?��3��M��W���c���i��-��0�q�d��$���f�#웙�]2v��n$��06C���tc5
��G�z!\�f��m�4��w)�N=E\e/!t��H�τ%���s.{ zN\����+��9�r�?��,��N�ާ��c�������å!6���:�A֭�+ '"b5��߱�hI$6U�:|'����\�������6d��i�> G.���4�m�	������ބu���`�	���3b�f�����*�Ь0�x��L-\�+����Y�����$��1�xj�X\��5�ے�U��W���c��x&p��W�-���A��-�r��Ib�������?�90�i�;5ge+����)��$���9,�?מA{� =���� QF׾Vb�^���h�U�xS�O���E����4�U�6��p���νˀ�}@u!�ޒ
.n����w�V��W,)=a�DJ��ϴ/5j6F�@�#�#iGe�l����/���weS
�LVD*mϧ�����2��$%�T���˥}d�z��g*�ӹ��|�e�Y_��a�wh }��[���\iq�