XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����sdÍW��o�����A��h� �:ϋGTt�@�Ƒ�[����Q/�?.��Uw���}T�[�v5�9��kDxH�H�.4���S�4�$>��BZ��q_k�Њ�W�1��*���>{�"��Xv<@��1�#L �#<W�ӕ<�)���5t�vT�Rr���B'��-V��{�m,��zojv�Gb���1a�]�k�J�����kk.��6�&����z�B��l��9�YD�|56�<��<8��v�B�����*1?i��.9IIw��T�^g��#�XVR�M��@��W̐bd������lIe�-ѯ���6�oǇ�Y���������@^AH~�9u�Όc��*ѣ�7��.�-�ž�v��q�n#3HE����>��[C�(R�%L����S�Z��T�zr���W��RY�����-���wQ�����<P5����׋�������ǁ�j��j/���E���x��F�0_,���E�+@��v�ֱ�&��#@���U	����̢t�r�1v�~�@��e{�~
�<�lŶ��(����.{г�����m���t�yH?c��"�EԒNS�ZC������H���MC��C�V�]���C� �~�1�̖�Jya��(7�L�}�E�����*Q��5�*4��m̦e��h��~��Cn��n*,��+�֩j��`����_�/=�T�f���f9�A^��'z�����;|�Ap2�Z�T;��������gXlxVHYEB    8e9e    1d40���1��jb�ʆlՠO�(B�g��~�PQ�`��0�'*��4CLU�V�pHL~���G7�!k�X�V�����)w���Z�l���&Nr:G�=�d�a�r�K�V��$��xdK�`&��زH���T���j m'�S�
dA�6ǘ�w� E��6WV7���s^q��S �d�߹]1�6`|.�b�gp��ǲ��uS2A�1TP���P%ƀ��j��K�w�N��}c��Z'�.�Z2� \G}�7	4�Ȟt!���&�F�f&�����������<l�Q��V���1;B��b���5w9�!ݎ�jG��ׁ;�P6<;aNP��1w'�������=8h7�t�'c�Aܚ�!�DC!ϣ����D���vw>*��125��g��4��'�&;dmT��0�*L�c`�ATU��B�̪���IϾ��R���)���,��K毓���D�_��P5����2��F�2��<l��^o��=3u�{�c�ϐ~��|��$WyR͑��H�$��ˡ[0��kފ�,�8��"�JAs�F��c.1���� _O.�O�C�a��N-%�,��نɣ	��Wp�#<Cn�JF%��T��,~�j6������4rpvԈ���8,�m��)�aE��">��Y���M��b�4
l��Z1ï��T���D����'��:��l�}���l�=���$�5Lߑ/�)��~SL;�b��EGZ����5�<a��L�Vc�� ��]:S�+j������G�b�K�X�=:sW4���̨���)��Ip�Ub�w��EYQ� *���p�J/�E�L�}Y pmc�7Iu���E.�Cg��ˁ�]Ԑ;�'�+�f���/;�t|���Z�
�tS�1�o��2t�J��T�İ`A��p�oHzAQB��Y���v�u¨�wZ5�cz�f&6�u�|�m@j�Sh�o�}�0}��؊�X|C�	��{��N��悥Áx���}��ޅ������D���jӓ�j�h!ϬiY^2�ώ��,�=B�&���+�Đ��t��y@��T
�\O%�������2�\'��kh>.���(Գ���v˽�ݨ^n���[3��d]�QO��>5_	�p�(�Ȍ��;K�TcG�m�rj�;���p��?)|��E��0�n,����'����to����A�ï$+��R85<�Ԭ<	3�]����X�v����<"hPT����¨i�;��bAk(�T�	� �/l� ۤ�?�n7� )����|&�i�0���I�)�cev7�2)t#��(ȗ�$ ���=k
�	�F������ �W 1�UŻ5�%���6�JL�8�Sʨ:�U�G�s0�Kӹ���c�igk���"^�^G�@Ն(�+ ���-%Z�ml5�*�߭�e$�}(?�ȍi�������rP	7/���W��mN+i�����B�3U]����-99��͕��jϲ������!���>@�ϮR-�6J�~�މ�qַR���[d�G7�1��ʛ	G����=�	jD���/5��n���~*��N(���љi'WÿU�x:rG��C̱N"3}2�p�6��YR����C* �s�m2�
R#ie�?up��.�T���0��P����u9�%�dp�r���v�m<��ʷLՁj�cS�O��L��n�E�4Ù<�g�����ݿ��[h�`�|}`�꬗��{�M��s�8H�c�fpפ�Q��/�N$��>�UG|j�7|�F[j��J�s|Jp��9�'��ȇ�8�#ݙ��c�#���>���f�1Ȣ���������x{�C�z�Ѕ�v�}UCn��̎�9 uWdBY���U���k�c�z<D2���ʩ�`t�C_r?��{P�
(���-���q�����6w�9�G���k'7��J��i��(x��F��6�Bp��΂�x܇�~s!)�:�M�扩�Ae��h�����z����	K��`����t>�I��1�)��|F�_��E	�!*부�����w�R��p��#LXp�7�|��7���5�d�������
ē=^m�V:���Ժ�90[�5�*�ʰ�حk��jFn����)�18:UZ$Ҧ�ޗ��f�B9��/�������1�	�h�*�8�bӂ���x ��0
xURxO���FR:Y4��Y|�q��"zd��ƵGD��u�H�S`֝��{�g�>%tv����Ϋbm\B��X-��x3 !\�=Q>�-N�}Y���a%Դ�Gٟ0�@�<#	����'������?�;�y���C��(�}I��s:�5�P��M��wH ��O�3��%�F"V,l���O3�5a��~�WK��Okf��� � �A���r�?j���<5M�Ð��L�t��#�U����9�9מル`Dk��ea�;��"4�/�GI��C\0|p���n(��W�	e����ғ~҈C����HD��46%�������7h��.N�;Z�o_���\�����{'�c�R�FB�hupI/��lp�2q��_U��H�Lԡ�x`_X�Įw
%x,���C[(n��D�ݡ������jn&��d�	�r�sxT�0���+���.�  -g�|G�#����g�l�L�Ϝ�ب��}`H�������]�	�N>�v��
��,&F��:�ej�Sv�x#h�����xcP�p�?�'���^Z�~*c���i;�M{�gб��k�KtN}/��M\IK��1H��XCP����cVQʅ ���Q�&w�$��>�-m>>�-�Y��!���*f�}&-���x��.����&<���88?:*��G)T�=��Ɲ"�-ߗ��v���z>�`�R���UmJ����C�ˉ��1�x��I��U��IV���/����@��OC&��_�n�A��^��OW�w4t_�j5?S�ٷ�*s��ى*��B7b�{�e��}��W>��<�0p1	i�$=���У� �������.v�x�XN/��	����o''���"&���VUL�wkvjږb�3��V�E�?èoR��
�{�zd�����q�Q~ڒ�l~'��>��h����J�n��:�e�4�nS�� :��.����rd�,ڽ*b�_j��1����;�i��0���ջ�J��0|�=e� ���Y���C+gmE,�	YAo���U�]@Y���.Մ�������7�59b����m.�6����9��\���(XZ�<)G�_n�|���D���[3n�e�Gj��˪vc��u|Q:P�G����Nɂ�	�:�\S�Pܚ�Ԫ��'W��]C���V��J>�v�x��*Y��o��<C"�wX�g���#A9o�ϟ�ҡ��,���ٜa�j�nnȵb��!�v�Uը:"�(�1o3�6���zN���V�p�_3ϯ��(��7I_���O)+5n�x�ŉʊ�����"?���/$ɵ'�nd��`"0�R��AU��6����>xM�&G���ȴJ8i�ΖoYEr�ӥt����c2;���>�t�q`��u���n��<����������E�x��gsO�ŝc4��НM�~(3�ɯ3�
�[����i�O����7(�s.u
ǩg�op,�6*˺�w�+��/��}���>��|#��`}07��C��#��Ȭ�A��n@*��Woᬄa�kؤ���*��5<�_����V�.���)ƕ]sf!���TZx���=>�M� ��VI����.;���=;tav�3�~gx�O��}�%΁]�O윑i;n��߾��h8���ª�K���R-�x����n���@=n�8�u��. B����;?�V��W��6z��PLy�d���;����;�8������1���!��G{L�O���X&c�*/����J�}G;M<�'��a�7��o����DO�}�&T[o���cP���a�(dN�^�hԧ�|9(���k埤};�r�`X�{���ӑ�<V��{0c�<Hw9��ғx� N4G�il�ד��_�5����3=��-�����j�3Q�Yc�,�9�_�q��DQ�Rg:��:|3.� ��[�%�1�����F!bPw�L��2燍�цy���( <��a�w�b��Z�K���t�P��������WǱ<6׬��HuGq3}.TG���H1}� $��9D!Q�DX��20�L��q�~�� ��R&9��F��9/�!��F2�Xp���Eσ�n�}�,h���1�C�w�h��$�l��q��a'��g�̀b���{?6�	���c�7ֺHf+)u�,��ƅd}'r/���?ȱ�լ#�)����h&0eK��K�8e1-c'���v�l�Ţ�e������%��X����z�WJ���'W���q�8h���B������A�����@]78��T�a�Z��JB�$�I�<\�Zl����ir:g\�3kA|�*���O�)��J0U�,ۤ���>n$�T�����+���=�cD�Jt()�>o������k.V�wr�%���>ڷ�=I���+�IKK�>�]�N!nxdg�����L�j���ȕ���7��[��|�vڝM���^Zx3�Y+l}Y�ee���� �R�ߒ�e��L�)ҙ07�����|Bu#����$��V�����@2&>���+�R�a����c�Gjq}v]5޹����0b�P^'�����Q�Cl����/&6\���f��3�h���)t|&�େ��X8�Pkʘ�ܼ�q���/ԍ�$��l�:�}'��r�$/a���qz���S6wJ������� ڥ�j�}3���!����%t	g��:>l=��pOGfQ�_�Q�Ax�M�{+eY�:�b_�	��h�e�jb9��28�m�n���+q���qj�̀`{��a[�ٳ��j�Gnr�d ��W1��9q�^�#B�7-����9q��B[���\����q�}|:V�b?���vЦ#
�Z�����P��6�᰹Aq����P���3�|�))x�x���Wɶ��6�)���&�`̵˔W�,{$�z�[���g�iUΟ��w"�����@q��L�J�p&#����Q�~�E=��ᵮ�-��k�&b	��)��t�q2�D3���/X$��kCE$c�!��W؊���BP�ݰ��l+��L��9����mEf���=e��D�"�d�C�䄰�5���5�SP�����#X&�� K�~��$���7ݓ�BI��G���S,������ ��b�;;i�,~P|\�63
�9R7띙|�Uh	������l�/Q߰<g��( ���&
%��ԴL�ғ	��M�/�'���7zR?�c��A",��6�J�%��d��0r�;�������l�{��fӛH!�_����j�2�d*����^�vd�|ԧ�?Yڄ{\�6��.T��� �xt#a�
�cm��s�A�DTo!��r���\��U��8������նsd��:�J䊕�&�+��Ҩ�73���{�k��H�:V�\���h��or(�r.��]w*�+���idQ&`��n��@�lR�p�������w$,g��X�j8��]�Y�$�n�~����H�$���7�Χ{�Z�Z���fl�ܱ/�����,`C�	�"Q�4�RP�R<���T�P�Y�h���DiUܩ�J��d���_+*6�� ȣm՚��Iެ��oo{no�8��;j��p:�U焞�qm�1`rZ�vFڔ����D���e�����{Q��w�\��Y�&5ԇ{oZ��茗ĒN�J��h�s��&a%�B����Oo��G�x�/��T�M=�C(r�-�4a#����h25Es���s�b�c��2+;�	�Ccm�E��z	�+I
����o�^����;j/��F�����oO���ٜ&(br���y�r�CL:�(��Ԇ�"K5��v΂	NK}g3�(������<O���Y+�aS��n�C�t���!b��LKY� ����i�����6J����� ��wx��V��M1i�X��HH{�ZޭE������+U�+y>̆��"�L�7��ee���4��9w/g�a
�Jp �+5���&Yfv��o������#a���/����_be�0b�W5p�Jl}�J��$�a�/�ʼ]�q�@jV��OΈIבֿ�ݪ#�u�r��v���e2�<�,C��(���Gx�T.���!:�7��2�mع�Ȑ,�S�oW:������y]~[b ��*�`}��v�r�TgnM�D�}���?�M����c�/�|����(ű�}��+nl�O�ۺ�����\�Y�q��[��+�kfy�=�~22��)��0�ܱ��x���Q�^�w���5�ћ�����������?���K��7Vt&I�R�F��yD����q��>}�fwf'�E��ɚ&�I	z���y��+U8U��_��}�qҔ���P����%%2�G��vթ*:8F��3�]���zC^����Fs�vAu�� �P�Ä�%��:w���� ׻d� ������!G+�?u^H�5��æ�8:E ��I�"߻�}�3��q�S=��\�l��
�$ҞjM����=�g�XC]��]��U#��&�J�6���~{Yè�8�q�K��Q6
MJ'�/*k:g��C��	�'D�M�����7��i�V6D�A��=��&_I]�SC�
׶�P��J�T���-���~V�o	��p ��
�nI!���@��A݀�mK���e�l�+X!��f��o6���=2�i��1���63A����)LÆ��b��_S�&P<j��&P�R�Sx�#�E�ͱ��|h+	��0��^G9�7��
��E6E
�xK1�����<�ܪ���/Q���۔4�E�.�J"~B�j��%C,5��9���V�#^�1��1����P��Z	8~RE@�F5��4�+�~�]�
Hg@V�iF	�ޕF@w�z�* �|*jQ��4J��bn����ay����4�����$�ئ�>�M�.�0{!�"��T�񳳓?!�M�$����,���͛e��*E�ˠ^b'���ʃ��H"�6�K"�\�kg���?,��XGe�f�i�6u�+��J����l�~�[��S^a���P(I���iU��Z���/�b� 4.�(�E��M6H�+�<%��S�i�%�&^��T �S�RP&�Vd������q鿊0�-��ʂ#͐X�]�1��w&�Le6��6���>��O����0����N��\?�����Hƞ����Ǐ�����Qm�C�d�j�ۧ�F�0���^��?��9�KdYؐ9��U�����1ٸ��+�b�}C֥��i3���v�%���Q�J�E��a�X~1���6�H-�C�E�f�(�oD���J���|