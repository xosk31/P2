XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��f]�F��7HK��N����l��d�ݥfr9מ}����ۏ@ބ�:'�s(� [��Sa��`��:����7�B\��AD�u������G�P�	ut\H��T���un�op+L�L Kh:|��[��iU<�D�Vc����Y32��Ӫ]Zw�����֐�y��~dv�\Gq��a�̮�X�f�P;h�1����M�*Q�]z��q
Ҭ���}�>V�hPYPl�(ڃ��p'xGfǵL�qceÀ�M=�G��Vdj'�S��v���MJ�g�z��N)���:�:ٚL}YM���u��_l}#Ɩ\.�dd�if�&3�������0�cE���*��Fr�OǍ.�0]���'�C�����0�͌����D�xDu���ӭ�zv���,�įZ�k$d��֨�`Vc4������
�@m��iZ����=��)��b��&|z��c&4��'ߡ*N�wr��qjϮ1�Da�(�(�~��ep��
�����"�&���D���MqTfN~.�ÔW�T�˪��	�T�A��e�~�wlxp�O�Ɉ�P~MW��/}ԫȗ{�>��P�����s��:o�=�� ��M��j�KeA��U*@�f��������="X�����O)�zqr�lYͳ�_Ω�̝CL���E`���C�V5��%=�G2RtZ�}:#�s@Q{-鋞��I�ʾS�Ƚ]�����+ٚ��i�Ӄ�bW^����2ĭ�M2CBψ>yz��k�(�?���5�B"7XlxVHYEB    1c45     950��m�?+a�0lFm� �Y�le���8
�Ê��9	Z��YR �î����n�Oɉ� ��
��%d3~G�����2Ȟ΀ѱ�'�i��/v`���e�����ȥZ�Lު�I��.ö��)���0"�usul3�{r���3°q�=�Km��,���+a�U0$؇ЯT����r�(��$ȴ��TO����ϱ|l��y��MD i9e��F�qQJ�s�Lt�?W�}���ܧ%4fr�I`�B1y3�3����5�zᇻ���ٱ*���P�3^ 8Ԃ�@A�2\��
�IX5�_G�BN��-�މ�k�%����������'��s��z�y s�h���?�[�A|~O,lQ7p �Ĳ܀r�ѯ��(�e���j��v���YD(sW��V\���	�.%x?�M�Ź���I��
�elz�U�WR�&�����5����2�
��S���65�m�Ƣǟ�ٹ��lol:���D`r�/���8Nhq��7b�H����yX������C���*�lU��r�t�<0�t�y8�U��Rp����#��V��<_�t�1ܾB���5*�x?��n��p���M�0��n��*��yh<�C���/�����Wr}|��١��j�Qy�߯�����@6���F��P�"�E_�M��8ZnS͊C#MIf^y;8*ƴ�&`��[�u@[�B5��ų��!��:ɘ�w<����f��V��C�j��VX����O�X���%�.U 7�d��;��8��'&��)�����u����X���M�r�[� <�ւ��S��_n���Hxc�� �Pȸ��lZs�z���K9�K�S`s�y/��뢝�y�p�k�DQ]���C�Αo���������k��0���N�1���;I[C�����v�}Ə�=�L��1
|�t�B��h��Zdep���x�͙cw�꜀l�C�E&���Kquu�����rE�:P�N�pY�i&��o�2�Iwbc��* �4Ab/'"��4����(a)H�"J�0��UA����/W�*�J�4'��K�][x�EӺ��8�-k8 ��w�lJ��i��B
{(��W�����p�a�ƭ\�w�f�_Z5��~�v��_~y� �Y\�@�6q�`�7uL�K㥈'>7�If �� ֡�_�ݢ��uOj��#&&��
��vmٖ�U<���7�c	H���C�d_�Y��`T10�N�O��r�;�;g�d��ܬNv zB_�[e<g*u2"��-rj��9 9�P��Q��0�9�)+��Vks��.�� ��73-T�[!C������6
$d,c[x^,܋!��DX�O�!��`�YS>Y�F,4dU�%�y,��5�� ;[T��քfb�:��Yɷ�*��ɒ�1#�8�e�ˮ����B��r����;j"1p��N�rL�������O&��G�|_�� ��^��.����Oy����rS)Zk>�瘝�9�� S�A=����٬]�Ĭ�n�~�H-<?�Ȑ�-�z�u#5/]��"$����(���9lѓKe��h��o�[i[\�,��3�.�(d�p�_m`���t7�qO���cK�M��� 5��E�L����G���ծ)�o����rU�X������;��[Þ�`gNt�������,C�
�Q��LӬ��%Hp�ev}�����;u�,�4��BZ�b��*y\���;��00�oy���ֻ{�(/c�2g���Er'�Y�����O�B�A�*�G�*��.��T��E ��e���m��ܳq�[x� \ �����c�y�{;b�MW<�Q�}���LAE?���7�=��?�G��'�tʛy�]	I�s���-�GX��h�+ ,��G0W>l��݋�2����tK����p��r�٬eiK���8{���9]�3$6C3=�_������]��1~����/��-bDQ79��JԶ���9$JB��=n��xۧd�%���t����?�K_�`�ɋ�Ϣ*ԆM�V�ep�+N6����>�d���c@��y(U��"��]Z�1�׈�oD,fb_"'"�y`�u�k9��
���j�I����V���/I�£0�t�w��B7�/W:%6tʫ�uN��MTO����j�~��%�s�RY�W�NF_\n&v5���	�6�LL(�2}�(�A����5�8�������hy�M'F+2��$&_0����gu@�]v
Z!�Ǵ�x�Kd�fJۖ���;������~L��"�����c��'i h�l���u�+Dl���p6��d/'����{��]��cw@#���A8�������;~�V�"����,�fy���N"�d�f�Z�2�}�����i^�@