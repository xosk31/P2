XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���r��@�	���rT�H�T�H�Wd���8yb20P�,䭮�wq�a?�C��������3�������[��ŐǇBUi]e(�z43����{�S�⤭#��x�_�o�"*��$x��2]d���sE�_o��Kĳ����:�e�!x��q�?�����Z7��A0�.�W��U�
�T��h��s�%���7]�K�/��W��ּz?�.8�I����LU�0X�d�o�qB&�+�)�ZS�{�C�]�fi��G�^�'[B��V��+��m���]:��t�͇ܫr�(�B�4>��\�W�gN#�z�C��Vp3Ô���˿��X�Ye� �z���������M GC�;�Þ8���l�ר��$��E6�Xko����T?p>�So9�\3U�v��B-���x ������I�,4k>�Bp�TDAX`���+>lo"3��j�i�wD?������9��ħc�%(K�ۄ{�kܚ�>Jw�D����ӌ��K���]u$ೇ������g�X���6�){D?)��n
�F�+�6�������l6��=�p_#��a/*��'���>M�o!;�߈ICZ��=n(
���+b�������������/�Ԝ�%Y�;�AM' ���O��b<��a��UΧZ靇r�"�G��r�Xh�}��5$���&���O�î����"#o鋃��X��o��jj�Ѵ�2����On�9�2&���@�YT��,��wjԆ�q��/�Y,W^"��J�����XlxVHYEB    fa00    2d70�w#�)�O7�K�z ����Yϻ��+f0�!1��3�.[�>zW��in�O�.�\��X��[��ج�0�S^j�]yG]�~��t����!��xv��i~�Ji
j�iF̌[�қ�-�)̀(��E�����S2y��G��R۰�Z4�?�� ������U�?�Q�C�����b ��<\���� ��M�RIGD���D]�����E��R���\��I��� �f�e��$he6ll�M���[ή��]�g��7���I��$	��G��('�2$u7.�yS��"� ?*<���I��]��u�"���'�o����*?������,�����������cZ���\T�3����.A�;��6�!'�?:���R=\+�f��;1��m�GI����YeY�x�My�Z�Ҵ���hw.�^�q�89rq[+cl�Fy��z.��D�<�����Jv�qqV�K� ������G���������Fr��e�yG���|o��)�ؤd�fc_[���P)��d$��K�y����w��jM��˟/�V�"�61��c6$Ql}ZL]ڬ�V�(��4t4�f�̶.�·3a�H,S������2�J"�j�f���Y ��J��	q�Gg5?m֧�5C5�S���2!�i�Yn�j�����v!�Ph�gF`TH;+�t�������t�hg�d�y�����ƌ@�&�%��ƀ������R�����B"@�]W:,-Ԝ2]#�<Ԯ��	���=,��������җt!���*yE6�HM��ׂ��C��1ᔝPg�B0�i�nu��*C 18�Xy���g&�n#"#p3�oG/����~�^5zB�y��T��uLQ<��]3�w)�CҐ[��&�q�r|zCV�1��+��O_�Z��))�o��cՁ4�.���r	B���·TP)�����G�C0ԩ��yf�<�W�\KT�G��H�x�G�FQ�Ō����]��[׵f��~A���S]���i��FK�K�l�O�D��⸋(
�ы�؇��ዂL�[��v8~f)�����_��;W�'@���GUQ�+h��9e���yX .���lzr����1�a���W����?���`o�d}�0Q�p��=�)���L\F^�B�5|4ȸEE���+*h:;�0H!��V�<�>~N6�Gy���?�,���@�}	�k�����x
�N\^�{d~�/���o�2$yJ�!��������I�7K���v�޺��0�X���jL����m��ϩ���V�����Y�8x�G
ֶ�C�5Je�A�}�l��Ƨ�����ム���I�qR��De����/"�?�P�u�'Q�n*y����Z���6��>�:T��^��y蔻�V��Z�M�����l2��R=f�i�&�B;Q�w�D��ˏ뗤Ln������Y���Z�-�aT~����A�(O�g����֎E�	�`F�J�-��
y��Q��j?�&�ٵm��w.�v�g0��=:������`ځƱ�ۥ���|�B����_�M"�d������j�u�e���^'��v�J�o۫�WB��yfOk�Rn��0���A�qTTS���.jv
���� ��V��D�8t�Y�*��k���)3�����Mk̵ҭ���UQ�G3ͦlb�|�e����f.��ܢ�4G8�rS��|��3�\��Pel�A�l+�`�-X���8=�\�B�������4�R����u`E���Ӌ�)	N�Ő]���}fs 
��q��	ғ��gy��I�Kk��d�cSZ� q��!��ќ,�E����E��7N�}j�=j=�ۿ䁞t�� �Pm�����{�[#y˩���o��73o�����~ͩ곘l��D,���0��J	������~Λ�M�����⃭��>�J�ѵ�=,o$J�p$?�i�ɗN���2%�������F�J-���W�!=d��d�8�n�W5���*K~��׈[Mb�2�1���7�]n*!��+��gw+LSf�
��O�f�X_�bq!�u�,�M�o�f�0^έr@�I��@�%�bt�y%������N_�ٮn��֙\u��=A��Ek&N:2ާ=c��/<T4���d�~�|�$��
�Q]m�Jv�/�}-զ6u2�Ԃ;��B?k�JYllZ���)��*|G7����#Mh��:��M�p[��� ��6H��'@����^�Zk��I[k�L�| �x�3���(� ��A�*k"��!>T��<L�eG��ʑp�;�����$/sRxD��!�|z����>�n�ep�Ҡ?p,{hC75�)�B�0�� �,Q��b����L,�H�w�>
=��j�i����%����B¤����x�
P�n��}�l�.����!j�g �@�3�wèݡǱ�5n?݃~V@6?2��yK+�dy���fBMH]G�6�r>��\W��[����6��DH��h��Xv*��0�%4L� ���U1�`9l��q���T�y�lSmO}��#�^T f8�u�qG+��k��4�`��X��ͭ��5��hN�&T��D�������}#�w/&���%�f6��hp5��kRKfa�u͠�$��.����P�.��^�=��BB%�{�%�Q(X�7|/M���$6L�JA[��a��0o�#ڨM��s"@�x��W�T .@	w.)�R��aɱ�87,��_�F)���o��]�D߷��$�_2����AyC�W���@��V2%Y�]��dR�ʢ�p��}�*s��븮��WXMm������u���e�Z��2Ӣ�P�B�3�6�+>�A�g���h(���[�P8�@^(W���wOǴr�����9��WoJ�����N��!ue�x����7��C��<�˵]��͙N�'��rB�.6���(��"զ��zX륎�+�7q3�����I� �H�4_�JZ��ܳ��nB�V^�w;���o��ἢ�Q� 5��6�T��E�{�G���`�@���D�Ϭ��U(����?3���\��3s�A��ӕxWb�LZ�����XV�3�_/�7d�>h���n�M��{�/82����>Bʚ�5�a\2Nb|6#��;�:u�Xpk0eT���P��q�l�̆�I��A��@�(">u\�j�S^����z���ŧ>�Y߰�>D����Gj��e��2u��
�I�6�;Q���dQ�<Uw��B��Fz/����P+4pnʦ�`��o1��j��=JW�1ĸ�Ϙ�����PO���&w�_ho%5���>�$�E�ܰ=����<E�wV/!�@M(�2.U���K%�.�1��u�g�@Ң�{�4ѳ8�hu-�m֦=�\�e~4��i�1��tt��x|�I��Ɲ~�'֜L��q�G:�^v�X��;N��A_h�S�Y���b&� ʪbݬ�l9P��Ψ��32��B�2C�1)�:=v��5_����?���)zC���lgx>���%C����S��!%MY1����N41[�r����E�qsf��D�t��+i}E�E�ص,i���	f�oo�g�M
��`� &[d��4K�W��9�s�r�:6[�Ҩ���숨���=<M)n�#��|����Zp�=&�~,��[�1��8S$��2��Jщ�Ku����ϲ9��G�<>ԉ5����cKu^�1��;$�sf~���Vy��o�z���B��Kb�j��*���3����I���A��"qn"�m	��PG4����k�,��|�I�'�q̓z}1�z%_cl��B�A�nC�^��`�>i	��
^�fX����Խ:���W�M8���������(��U�w*��ɒ3���6cR����p6���q}���n�Ε[���.*�-�Q�1��}���qg2//iR�Gv��,d�^E�]��	�?�=זs 9���H��$Ώ�	�DJ7�\�z(����JȺ��䃬m���fa�>�>��1e�9�kY�$m��+vs�X�Fs �W�t�<�^C�)(uD���+N�fx�ET���h�m����w�*܇��![%�j��m�C��h>�C2ذ$sLk����<��L�AU`5�V<l��ZTX�C�KҏwE�m6��uh%Y�T�.�{�NQJ���O5��4�c��1S��D1T����U�Zc�DV2ε`5�Ҳf/t�C���r�>�9��1�	��L��\a�É�v	��a�H)k&Q[$4�_����D�^]�stE�2�� |���4�.�df�N�:WpB�*�5.ߓ"r�fN }�s��&:��7�|G�ͮ�x��
3��X���E""�>Q���*ʃ8�V-i��X@��2�kS{g/���5
J�k��fJ?A�U:1T���6=C�^M�鷺A;	�z��c�q�{�kO6u`�(7�p��L+�v�U���}��	="+��GMul�rP�x?'�=:���W�!��9���>6M7�*,\�t��,U`6H����th�vR��h*v峢Î�x	���-�CEὫ��l\�,&R�y�t6���9[���ƿ��#�Kغ?�����n8ږG��-�XK`Y��fS?�A$�_!�-{s�jg	YV�8
2L~���6`�W ���k��a�*[��ݓ����A|�J�����Q�~������!n|��s{�u�.Q���ǘv,cŪ���J��h�!�v�Ưw�{��1�J���C ��;40���T���EGw��%X��"��J��	��<E~��e�yy�A�a�5!cz�  
�͘򊑁SQC�H�&�[Rz��Ja*1KҘ�`6L<4\ߝ��@@�ꏶ�a:f�_Q��_a ;t}�F�x|c9��ڂh,�4��v�:��)>cܜ�D��+И�v��4ڟ�f]ؾF�����7�d7�L �mY�`�}tŬ�J���n0O�������+��1�L��\��B��q)��D�${Wއ�|-����C��n�'g5�S�W.�<ږR��dS_%���a���;xK�#��?R�d���q�IEÅ/VI�V�Gwa� ԓ����I�[�W9d��D� a�jA�1��N������ S2	e/r{m�X�����q�����4�$�B��2A$�č��ݷܡ��s�O��C��Ҁ8�s��P/��	�s\�1�CT���ޞ&,���mC����ut�� �h\l��}�JH��R��n�UOVD:V�����s?�X��B�ʕV����{���4�z'�7j)�?���'�����
Ƹbޠ����V�tr(i�[D��=��� e�6�� �mgTs��2��T2/��*�e�*}��[ZB+N2��h�Z͂@��3H���*��+�z6���Us�Y���V��ɝ`�]&�)ᓁ����f�򁀽��"�^�Ƨ��3�l��* wd�'O_?34-<�}��`8h����QJ����$������`!m��9�uSY��H��lV	P�2��3_��_ǟ�DU �d%�u����#$@Ty��JvNK�6!���Y�g�W9�	a}�>Cn�Y9D��K�{o�:�x��[U�l4�Q�����񓩜�K�AL����NFj��T��K1���A���[�=�`�!6M���ou��8�5��d,$ޤZGt��-�"����S���ŇJD�G��:�fd��Ү���ͺy0�Vkn8Yc���z�@���=�7�U� rI�
e0"��&�1���Vo�r��`*���#�X t�gW�!�R��<�eADB���4��+n>fOV\���B#mc�+I%���d��cSܮ�h���yj��E6����"�����g.����x�<��y26�<:TC����45�Cށ)%*�$MS��O�N;��:��<�ٽ������T�X5���@6��H>�33�5[i&�Z�v������a�S#^�n�R�rCR��+�1-j���:�h�4;�htKݥ��B��L��lQ>{�=�l��j�J�R�B�����!���^awZe����c%g,�	�?��_�s��_n���t�\�8�b:\7q���)G�0\]U�泊�g�GZ�7�89�s\F��E�hd����^�o2(Q)���m�iM�D�M�V���!8&ۉ�%չim�8y��҇x��*l���ie��f���rOl�.k��PЊ�t���P-�Q�ae���+�@�Pb��Aj��� WbbF��w����U���襋YD(sdJ�?YGM��%�߃e]�7���җ�`��;I���j�����z��,�bR& �\z�BvT�<{
�RX(�)�y��9�G��'NPN�<p���ۉ�j�X��wM`l���~�{�A^,��dF�F��~�Q�5Ӧ���^b$꬐?��gi?(�av��eG�Y���uB܉Jx�e5u&��ZU4Rq$ov��ф5�~�8��l�"�硌Q��T��n�c���%�N̾d�5r� .��~0�)���-��YݶaD�}�R	�f�$�a?芦J�ӵF�[���(z�@}[X=��W��ƒ4�)G��K`4�Xn�@�9";>�l�g+}�ثǕ+	I cpn��ǃ�!�W0��D [��
Pc�v��ˑ�L��pAY�	��.�b�Ǿ`-�=��io���\9¦y����k�c����h�I~�Y�M�'��0�<��(oaz<�|�3Mx����=&��B���iX������/�J�;�s���<#V[��6{I��U�Mub���"�8f�PJ>��~,d�?����?��&��s
�����Ŋ�xW�����
��
�a�҄l}Sg�`˭��"����i��2KF�Ͳl]�KQ%�q6ޔ�/Ό�EC�T�<���{IQM[�U�RNFh%�L��"�������K��C/��@�91��.Ȋ3��)<p'��a�k�|ܓg�q��?̏��������5��F��K��`�{���3r��&�l�t!�;s,n����&����2ƊN��h!
U?O��z���WjUg&U%���M3�>�*E#ztʾ�2�Muz�f�J�O6�qݻ���xV!����C���YXHz�&沔m?)�#C�/�X��,��YPh���+���tMa�ɼ�=S�㛝�f���Z��;��pZ�>'b�L�x�'=�-��s[,��j�$��	ie�V�$�y(����מ�y���x�o��>~t����f>���.+���1k�c�;c�y_X���hqc�@�ςn�e�R�Z��v�2rF�J��J	et!�ώ4iE:�=�D	x����`�i����x~��d��%�	�0��/:D�t50zI�OY�iyF��~���o��]���2���#cI/�`s�z׵4Cm�Ju�m(e"+Х��9� 2�����[��3j2��}yd0��h2�ܣ)�x.P;����wQV�ISh�+�Z��n��;�/h���Tne�A�V�W*�_��쾘o��A�L}r�3rU1���8��Q%��V�c^: ?�4�����
�x���y�%E��o4�~2���y͇B���q�9?��j������J�#L��Q�_��޴e�:�CW ��i|�ot��1H��֠*$���U7y(< ���'�W\�"�xA��<t��ݲ��*��� ��W���L/0���dY'u�jq�EǶ��M_=Iw�)���/j�P�cJa���GL̺�*,���mJ}�3ٴv���Y�F�8��W�`�����ffl���1�����pj�*��"e��������^o8�A���4o�*}������k�=?�9����ܜ��ܘ	ZvD��w��
�d�;:h���6�����c��I@���!��|:��@�q@ƽ",9TV#�о��v6ݮ�%���|���o�T:�5#��X2 #A�3Q�����E�ÏE�3���]��*��]!h=����؃�dh�sz$��̲\����Ţ7����xƞ���
�7>_�Ĉ苇����R����-�펷Jc1����/϶�>�GL�>p@�x䜶s�5��yf���+\+6�L�l��BR�O)�fH���)oxx_�B���֖����#=�oN�8;�8}�eOA􄋰��
8�\��kd,����d,U��sk�E�����9V�b��:l�b��OpQ6���1�W^�,>H�It����[?�ao�'"�d��9&�*O	J�v�U& �� ���LM��}���g�y��Y���ǜ���&D�˴%wG�UZ���W]��]�Ah�:�{I'|߄����f��̙2(,K3�CS�F��I8*�<2ռVYW���XG��M����$���|I������cꕺ�����]$#7B!��~Sה���|���()HQO[g[�X0��S)���&mdń�([VG��t�<� �7b�]~���x�uxB�,i'a|AHL���_�ꎽ݊�=���ݍ�V44M��Gh��j����D�T��,��(���8���"-|��:^K�e�HH����Mh�IV΂�� -�W���h��@�����sQj����#ê�/pw�v���]�P�rʩ,Nk����뺫{��N�r��UC��?������5C\�b* �2�q�hzХ�	ud`���_���G%HK�g�d�:F�a|t�������1�vYr���-��w�t���wu�paZ�yf��ݝ��0�!\ �`�1u崏)���-���tx��V�Z����򫓓��9q�XT�����GU�X�l�0�\��Ce��ȝs09��'�Sjpjּ�J{#w���^�j��bE6i�<�(dH�3���GYT;ȞĚjǀ�5�Nb�,��'�wY��p�[_3 mi���R}&��I���?�m�ʠ�?+�1~n��a,���
����\���uC��t5Rpw-��6����h4�����6Ϸ��b�����O��� 3_m�G��9![F���<����e=o����%��Kĳ���}~�����>�-�:��d�D���u�cf>�.����[�]`�]�V��H4�k2G�A��V��u���Q.��;���-q����e_�ay2���Y�B����dʻ��/�D��8/D�l����׷\�c�Jؗ�l�p��������%�jr��z�T 7�&��T5>�t�IgюV��I�VI_���0���\�B|+wH��*-�a>��V��!&M���I_5�!�(&�����0k\�Ы���&�R��[w6�h��\>p݄����Ab��-yԔ���ҁe�ͺ��	m2���&�sP�l4N�A�07�<oe$π����<�0-;�X)���\Z3S�r�ש5Х9��U\�f��e�Mʇ�6#�>����
���to^ V�R7��M�9mX}}��Z�C��<Lcwi��=u�#b���ᴀP?�^��hdE���ɖB�@���;�u�wS9`B�{�G����ugJ�i�}��r�K��ĕ�$̻�h׃%l\��"��v�o�zɟɜB��Isa�� �
�w�"0���ǃ��ZKf�۰�)��e���JH�B��>��̮���>0�N��Ө$�_�+���}�*�{�#��0P��k��3�)_�xj�6�P�t�U�#M�7Y�+e�pJ���v�NOrU�O���bL�/3f�6��ѹk�X���ܲ�sG�4�,��l2���ba�A�`J�b�H�(�D��P*��kD�f@B�"z@`�M�H�~R��|Z6����X�J��x�=��|:� 0��L2�5#)��)���Qɦ�s[(��q):F�ٜm�"��7�/��o*h��pH!R�2�s:К��%�:E�+��^�@�	]w����)�� ��xm��m�}
�]��P@���E4n0��[0ϵ���S!�t��3&pϴ�W�f�æuՉ�fEۨ��Q.�x#рɁ�K��������� ���0 �b�:��~W�N)2V�#�b�"
5�˅&�{od�rJh�>�]E���A�����訶�W�(�*GΊ�%N\�cj��<���yU�6�I�:�����qǗ��!�Z7lyN:�FH~����E��R�8�0������=e��te��w_��ȫ�5(E�^���OwN�����W�#y�G���8��w�KZX,�)=���԰�M]~ajȋ�tr�o����烒��ۼp47�Vq��RP�,Di�&���zϫ]#�F�U0�=��S�i̕�50@h�ಹ�˗,�X�l���nH�B�
�z�z�n�g�����L�쮈�/�JF��ϴ���)�ڦ�r~��'��}�P�l��D��[�"%�4��w���G9ƌ���2@�ϗ���9�䮽�+ݽY5#{,�
���9���8�@uB."Fr�ówr{ژ�(8Ѳ��N���=�87���ݰ�M$�rdU�Ĝ4�!�_,*"���]�T8�#�/��Qz]9"ť�$�HD�o�\��le���bO�,B��\���t�yT�[ &.L�j�N]�|2տc1l ڃ���pQLt�� =HR�P� ��@��y��� o�~���� /Y�|�g�:�O�quМpC��
>�x/�pJF,3'�"��>�'}�2[�(p'���
�C6����$R���tB_f�n���ᶳT�dTP���d�5湶�%��bw& !ؼ�O�+��[�����Y.4t�%����j����d���+��.Ĳ����V���+�]�	#���JQ���Z�m�]�D{�F������h�HG5�`bp�|�~�c�)�<r���,4vJ�9���,�8�#���#��ǪU�N��G� _�*��`D���[��¨qf�����\��>�'C|���}�=n�1
r�3�R+��&��s�v�
C14>����-�j����*�������l���6�13>�v��me뷥�5�)�S�K|�D'U�Eh\�O���i�f�ѸJM
D�A��M�����x�.���x�Q�VR���.�whC��"i�b�^u<�>{hH)u#'���-�{h�縫B��C�I�rL������O^�ķ3\�V@
�ZУ�u;.�L�F�T��h����D�?���=j�^���,���}���o�-�_"�����*�g�MR��|X6'zx>���K�,�y4���9`m:�3+SHaP
�%�Pq����]��f���U�H��D��;͟䤆�i+�t5�U�|+D�+�8�^`	��W��&����
״�w�=g�3�H1�{�j}9&�Ӡ�R������g��9sq�j���H~�)_��Ӧ���Ŝk���xFu?������\�Dټ��agf�Öza���xѰ7ؕܬ�u�s5�
�\�{7�k��|�[���Tg��M�4�Kܵ2̖�U�V٣�рQc��yސ�Q�|�����M@Z����3��J �hR����)�@NW�+�ͷp��v.S?���Oc�����]���@���׫�	ϲ��&���+1j:V3��C,]7����	93�'����l7���K>5|���XlxVHYEB    5902     f20����A90�Fӿ�,%F/�*̫y.Sy�p�i��z�T�|�:/(�����=&�'�?���Yn���[��a��7�E�'�.� �-�Ry�2F���o�R�P�ַM�mp���^R�`<���F���BwY�*�I�S`c�qT��ƥ�km�Ŕ�
�Olg�U�X�A�Ib
ꃣ3!���eO·G��k��uFA	�,P�}�a�G�zvyj��7��i�y���'����v�=R(TQ�w=4�Ո6i��BN6W�A�;��&\�� !h�y8t�8�Ʃ!��8�>|�N�ŭ//�#�E�*SJ�l�١�0'mAC|�Si��4�j�v�E�"ߞ��gZ�/7��Î���JD�5�������[�rL�}�M�62�_���^�R�Լ�O\<�r�xA~qq�4��a`��G�C����֕'�X$4��� /C�XY����	 �U׬�<V�X~�R�8����%�=]A��6�ЖQ��)�����G�0��k�48u�u�A������N51��C���K�줳Wc��X`��?�%�{��� P�a�i��s��*������Զ~��<c�!���vM_��g4�̮3�
P����<�\�����0�����W◻x���Q���G(I;)��
��jv�~F�(*�ǓyG��nD��nZ��Xk	o�Nŵ��w�F����0�|Z�@A	[L�p����V���9g�<"�~����"��d�"'�8��M��9\��ܱ��3��w"�(ǜ�����XL��)�.�10 ��;�x��ٞ����'_	]^)]��o
S�2pW�&xh���B�}��Tt��U�ɍJ�Wһ�))	���1`(��/���� BTǊ�U�G�1�>���t�Z����	^����d������z/_]_?'��r�΄`y��R�bK�����{^�)�8O:̖����;|�8p7�b�h�:������MT�����w�a�\	�z
�zw*0zof3H��+sz����pNF�������C�����Z�\�5��{�xRX���/u�f�1 �Üx1ϫ8{T��J%�Z����Xi	���k��Rl��%�lԤ���D�zޞ��*��2�YXh9i9�zf�^y{�ٝ�Ɇ���@��ش�%0Ga�Q37��(��%�N���� �y�e��P�V.'J��,�o����*f	��:'C$m�\���u�3�o���7�̠)��<��ہP��U��Ea���i.��b1ݡ�<xݕ�c�v���v�������e_���O�<Οdb Y�^O��߳{e2���#��F¢�b�b{5|}@Q���V�%�kt�8��aMo���0J*T����TY��9�)g"l��n�\B!3�>⫘���OwC%�G|u�):f��'��y��FIY���Z�� ����ޣt���[�D��BQD���x�FGV���ewL�JFͯ
W%��|�\��H˶)�p�@�Ή2��[g6%�8�N���JE��]8����{�-G�xik ��A�w���&�S�z;ض�f�h��Ԡ�3�B�pR>oʖi?��W�y�6f�HS2����ʾZ���xF�[3�O���{9Zz�:����f�S�R1f��Դ��2�Z���$�q-1� ����UL����g���?�YDsq�?Il��^
q���^�aӮn��Q׫1����l^�B��!W�Eos�d�Үt�ݖ�R�{7� �@�S`K�3�x=l~�pp&_Bu�!b�-ޑ5.X�ƫ4��e��ֶ%ᱵ���S����<j~{�O��s�=XMY�!$pEP�HLƈ�=E���E����'��C-1��C�b'�Xq2�i���ײSJ��òt�T&�O��ݗ���$�Z�k�HA��mu}���@�
�P9eW��+�ZM���P�qI{(2���pN�1�|�!���%���<Q��2k9�;T	�f��b0���0q�4pfA.�}��Lt�.�c�ݺ�^�r��a�M (�H�!uCTiC����S���%E�ԩa��p����s:z?W5Y%�&["-^�f�~��fior�=��� CI�f����3�,"<q���D�ٟ8��T<?�O��
���`�b
����X �B�ƫ|W����P��0�N_����nBƂ#��9s��Yc�G|� �sA_�4��z?�Z�7��oWғ���;6�g���2L�l8�� �ynOX�� 5ږ�/�ѡU�#�p9�JΞ
��vK�.~�*(��[ ���J3�r樦aA��v1���H ��Oօ���G��/{
(������&�Ni�-09���?ޭ��c���B��Za�yo9o��}���a�4�ᒧ����lF�v!�cX3K���k�w��ZP�bE<9��r�����8&�H:�7�Φa�Z3���m9�����K>f����˧?8�-�`Qs���%PK��Q�6�����հ�[�>��2c����6 ¥$>����Ì��rs:J����ѫo���~��>��=�d �y���������!��|\^>��d��꯼��L��-�$$s���.sS�#���N�'9��?m"�戝؋y��o�ʆIP��[�N3�u�>���I�:j���m��F�˼Z�%�)�Q�I�O���;��c���MX�gPu�*��ǁ�8�Y؛熚-���|yB�m=��á��"d�kq�]��7S��>����d���남�FC>9�0<�e��P�Vt׸���{��� 6{���#@`y��׵�3�v�Q�h��Q�y��\^�rI�MC�$���R�iV� �x%f�&�Ă/�����v�/�c8����[A�#�j��_,��g�̼�D��ɢ�˭��l��h RT����5�.%jH�v��!�d������rh����M�s#����mJ"ſ����A�.X�W�2~��i�,1"��K@!�i��@JҰ��뗗��M������
���o=Gl��oZcS)���Z]��������ll�i���G�\%�'��+��_��zE��^;�T��`�9���iZ%~��K���$[QD���dlp)i�b��R3F�?*�dr���Z ��`���_w�P�vk7=�1i��X�}�a���&�`��k�D=O=��t-��<h���^'��h��FOx��$��T�f�=���1+�>P��L��ڟ��+��`�=�A����y%�j�<׸�$r=�w�{Y?�pCnГ��i�Nv�vɛ����^��`�[��{�.s�`�r�'�\��j��"�����h�|��dDg	�B�S��5Ν�m]�z
W�
F ��W��sv�WX�H(v7JƋ��Q�����t�����י��i!�pq.�Vp L� ���B�L<�������g`�b�A�+�y�m�"�W��y~�*�?�T#LT+��)i>Us��˂5g�*p���+�Z�B�M��J쐟)�$��C2��-~'�롖n�e�a�-N��e���:e��x�(Yᛠ� ��v�(7��7?
���~��YWczb��b���6�S��<��?����`����t��1bm��V�����5E�Ge��F*���/���O�	̩QClX0��%^t�b�t[[��^*@}��CЁ�x����B�p�k�N���A�E�$�n��{�z���P��oZ'� ̕�zn8��#Ȯ�4�]h��Cof��P�J�gP��?E_��{��=V֠�lC�9��5��L=�V ��o�B���o۔����݁a������c�F���p�.n�:�*r�8k`���0@O�