XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���@7,pP�B�e��1A�����+$ܚ� �M�OFR��$}�˶�`�=7d��y�"��0�,�uÐ��OG/�r ����I���	��M
�R��.��ӐrҺ�ʡ�������t�8���F�ls�v�
@ԭ<�U�a�j��.�/��I��<�< ��eW˒#2{Z�!�f�p��a����p����ؘ���8�,�{%m9Bxv:��'���p��2LG�7�"`N>ڂ�6V�����f����j)뽄I�r�82�M�����S�Ԥ��6g3R.�2=^\�g4��k5���A�#=�i�)�~��G*�ڒ#�����)�b
�&#͐��4#�xn|KNK۲��K�ާ	K1��s����\+g(��i��H�Ť�Ϭb�PO��b\���j��z[��>�&�yc�Aq2��n6S�Nv�������B�#�[9�)��	�Lsκ��QN(G�~A��}��W�	��C�9����$�DEsH|'n�O~\�\Vj�C�1	 �P��Qm�E!���|����b�kÜ�KJSd�S�C> f^�S��j8�7h��\��ƺ ��k1p#�ց*�׫pg��R���Yk�(��梅+���;G�L�@!'��	�2�ګ�OM��������k�N��J�q"��!\��67��S��X�s���_�~� .�+�pB ��oiz9!��g�?-�����r���+
}�������)���f n��s5ߊ�3���<%�H���R��`�_e�e]��j��nXlxVHYEB    1802     830(f��? �Ws�ͱ5����{~��lB�^Ƙ��S�ղBi&����Է���'%���H�ve!���m�Q�lt��!E�|R�X��*W-C�����IaLb�xb!��4��x}��dg0lч���#t����jdL/�U�o?2��#�	��.�a���3�(J	I��i�H(���W�븧a+".�T��?�2EK��C|�C�a"ޯ�0��k@�W�����*�����+5�ŝ��C�ތ���yk�e���OP�,"P���5.���������Kń9���M>,�}H��=~��ΒrCԋ�v�U���P۪���D�,1��>�d�_%�5�ߤ���zs����qWu�aϗ�X�OyP�c�;��G���I���1��	��4ֺIr������ͷ%G֯�J3O*rU�.���u�}�w߄���
¦�Z�R��i�Wྨ�O�W�C�{ ��k䙲���?����igҎ���I��u�����j4t��8!��O�I�<��"g%G׃���8A�f�#!U@:�F[�4�j����ע3�x8��F-��y�dtY���Ї8��2�a^����a7��-&~5	���X]��KD+��K�Ⱥn�5
�=��^۰�0�r*E�_�}�݉3��޳��d����f��k�cG� ��|?7�ÌF:6�#�S�<��ԷFma���Y=*c6�D�7X��/w4��	���M\ ��O�i`�+K����1��n?� {���V���ݶȉ����y��U��;m�tC����4�7�!DED�T�Τ[��wm�&������~53~���xrxqM��oI㢌K >����1��φe9��T�a�`���2'�N�h3��P ��xs��O�nF��|e6*���Z�����su����T鿲��d��S@3��D��K?�~w�f��s�k	=95��+C4�J��j�Ю���h�X'��ʛ�z{TY�d��Gp�5�O�o���BR�v�pZ��}X\�[V$�
2��?+��qx�	b��`G�L��EX����l� }�.�?�
 ����U��X�䊁��"���+��zD�vǖ��	�A�HW8h���c�$�N����D�&iUjB
|�Y�/��^���Z��u�><T�Գ�..� ��S�*dA���a�6��o��-�R�:����.^�����Y�HIxx ���E���!R���W%��|b3�SS.�����{{��t�PV�cF�ܝ�\�OC�q�B� O
zA�����Y��a�v�z�?[�ћǠv�Q��t�¹�������>�9����a�o��f%7�q`%��_�ʣO�6K��S�\ۦ.}K�Ew�z��L�$]ꌨ;�reV��`�*7�k��R\�p6֣���1�Am9do/��㻺*:���٢P�j{�B-�o�/.�B��_\�����sZ?񇡅�������[����k|���q�~ڔ-�+,y�0߯��K���W�� �͑ʺ�W�+���K
Ԣ&O|��nɁ[Jx��6�~��`�o��W0z+�yϝ9(ԟ��|K��8;����t+�x���@K��L��Pɍ��9/����%g��$47`�Н`��BŞ��Z�2ڻ��+8e����BG�9�A^C��IX��S�l+a,Q�w��S�:Z5Z��rע]��>��$��e���g��д8��(�К�R�?7,qՂv�[�Eή8�J��l����� &��ˢ&[�����}�:�*��*�t��]��fI@M������"�0F��q����Y��ly$%s7�:Q�F����dz|��}�4@'J WC%k�R������s��Y�v��ۺ�^��7F5-Dݧ������
�$d��.��zt�=49	�����'(N5�Bҙ��}�*5L���
�&O�v	s���_�\�IQ("�=_�jW��OQH��Co3�+�idfx��`a@��a,��F�F'%{wZf�������Y�t�Z¦�]���O���y��ڥ�6��J��_��W�s|՞Bַ�Sy
R��E0L��eou��ᩐ�{ҹ|�����>^G