XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����uh���5�,��N�2F���c�R*ʧ�i�8a���0�4�+aR�/h E���*�%��,L{>�,	��~����jx,�_οsi �{��4���M�?�7�;��}��Qx7I�Jv��ޘ�h2�i�J��ߴNӳ����Ki fG��A΅���QPF�����[t�>�>L���>�Q73қ�&G+s�[�g��g��\W\n�>x���_ʷ*Z,(��4�hS�r�/���NȒS�aC��
�\�Q<�I��9����\l�L�a镁�|%��n��#�T��e��p=�g�1)�#~|��cn�6⭮�s����n�$l15�J��W�_�e������읊=��0%�a�/;M���mi�� �Dr����+mԀ(�SΨ	�Ce��T?4����iY{�C�0��u<��٠7�*�Y�|Dm����s�B6C\i�3L�����$@2�Q�z���g�S-b|�T��y������(�W�q��/��-�ՙݎd�b)"�T_r$[d�=�gք���-�R�@���J�>�{�@��c=.N���I��BՍ��K�ї��'-����oY�>,GŲ�ą�ɉ�^$%�`\��Zc���'�KH8��̊��G�?����: X'��vD�י��,n�b�ӝ����i���/�dq�ma�
ض��B�I���PL��E6�'���N�7�31xb�@���������D;��h����t����ַF�}�<��W�om#�c�(�S:�r��XlxVHYEB    fa00    2910� ���Į�抛����_.��Sɳ��|����;��:�4
�[Nk�)r�4�m;�M;��yأ�#��d�`�5ݯl���,XL�/-\�S��� �3F$���Zk/���b|[r$��%�[_��dدLԥA(�T�@=���^b.A��&�i2���9���C }�.�Y���B�����������t�Q2+�R��f�Ѯ�E�Q+Y�Z�C#Q�Rr4����s��������BF��9%=��#�ޜ�C ���� ����J��Vȟ_��JĪ�P!���MV�L�8 ��Q��[b���� m���l�0��l�,"jI���޲]���J�K��ǀ	�7�|�;:ZgX�?8}��A][��g����?�h#]ִͱ�����k� �]�r�U�tƤ�\��N\��^!"Њ%�ؒ^�{��Q+�[E�j���ӫ��6�'Y�u=���oqԸ_�&?L=Bs+3,��^�o��E��� Bl�`G�7h'H�����6�C$�&�"J���ѭމ��l�Zؿ%�fH3��e=��pG`y;��oY�E��űkW�O���1�;^dg�Q��{�����Y���G�,r�� )7��~Π,���E��fo��	�@TA�
�/�R�k�W��9n��4�	k ������S��w�Ϝ�`d��ܭ��g ��mð��$��D,����Ji�Lw"���G��g�R �yR?Qܴ5��o5ӿ���#W��fP���}L�6�Q����8A���<�����~�z���zr��Q ��*EH��l�O��o�������x�\�A� b����H5z� `���;�'N�z�P_X�kW��xij�8�k4Q��e��{o�饲�B��ֱ���N��l��51���θ*�@�� ��"��C�+��`�va��j,��W����茽l������֮_�ňB
�P?��E/���[ٕ:�K�vFI%�N�����oǗ��3�w+$�^#8�T@�V3��
�(��ۥ���H,��"O������h�����1�)H��^A���Ͳ�ėPv���D弑!L��P]��c
o���M5��6�<�SZw}�&��%�V�a9tH*χ�5D�K騒��7r���;S�M�mE$�J�٭b��jZ�s��Ɉ��qo�{j���K0�i~�<F�g�{���I�3߱|n뙭e�f1��K�ّcC�G-��u��ya�@F����Xع���rE�"=���qx��L�1K����ss��A���
�Fm|�O�ˬ�������Q~�%���:�
����z���`&�/�xHb�4��7��?4I�;�4��L�R�5^�ppXF�<لA��l���F6~��[���#Ұ\z�sܠO%<���DX�M��}�z����;�`�%#�,6}�p��5m�f�B�Gp$�	�p=7ER��7 ��Rs�z%D8���+a'�1Ҿm�c�ZM1�l�`Q���E��C���Ϩ�6ޔ��3�<�g��[���<���fKS[z������e��x\Fޫl�$d@���U�б�+�ش�m+V�p׺�zz��=ږ�c5�k���}1�>/CϦ޿~�!�k��ՙ��S�gg��5�4z��(.GO�13��Y�=}�������!��h�9 T�����ԉ�G�&Y�{����D���y�G�D������/^h����R��C�l�0i]!�<S�!����w�U}k�`�[	N)�>z���ӯ��bF�l�j� j�l��z�>|���U��\�g��J3#	v�J]�V�
̼��?���F�����m�f����j\�������{G ��@r�.��1�ֶ��B"��F{D�T"�����C��7Գ�-�J�H87N�e�Ɋ����`Qm�l���o���Oxd�U>�V��Ӿ����"I�x}pq�"F)�$� ������B2�]_d��l��_�	c�(����y�d}ck`����q CKf
�wJ�a]8X#]i���2�?^��Te�[��������ΨB˺���#����6���N;�|Ճ5&��6�}i�V1+������~��f��������`QX����W�c1D H� �6��/��RsQ�X��#Z�c��k�BkÆ���W�WM]��v)�B�(�sQ�m�w�Q� �d���	�Mzy� I��߆~nq~����I}��I�F-�>���8�G��A]�%~��N���"Lk��.9�!�����V`��m�;����L�2z�
��llo�1Q$�Qm�?8����⚕V�Cy]�c��e6=&�~H~+}76�xղ��h��)�D��Ei"��k)u5U��3$���j��� �M�`0��\	�ϻ�5�.M�qv��Vd��~c'�{�L��Q�ϕ%\±�Z�q��wͶn�V�8.8�r]@T��~���.�oP/���U;��9��;�F��%�/dfE�SZ`<1w�*���abD�~R�A�N����DQN��K>�!�3zK�u�U�t.�?Z�á�	g�_�e�D�i��U��V*T�rl�=H�S
��a�g������֚�;����Rb��b���޳�����7��1��=0x��������탗s��>��j�<���a��25b؞����0@����v�;9Իɾ�^����T�Fq������w]ü�1�-k�L��_���_K��-	�.�T�(��ч[)���!$��q�n]���J��kdtW:�rxzc�I�}��h���������c38����1PtJ�O�_���ӖX�l-������E8a����s��$<��%�����;��i]�W݋u3-E�7#?��u �N�a49~�m���}5����d��'�)-��~٘����͟�qd�-EY���J�z���d;ѱ�����h����[B=�ƙ����Y΢u����e�D0�w_��ı� ����fMW��1�b���i�Ғ��P���S�n�dsh?�'#~.��s���}�灪I���i5ן���TP}Q��H+G��y����:Am���'�֢�'M�8��
h/;��h�'�n �Ip��1Li�}Ӂ4,^|��Z�;[��=RG�Q� �m��w�I���萣���߈%�_u�&�ɦ��ɴ��<��_9����a�(�-�� �j��m�TH�Ja'�3�t��՞�󥎦�֐��|I�)7|�%2Y�=��k;�&����@C�W�>�R\�4If§t��
��ߵ��EʭX� ���W�r��QՃD��qC��
F�b9ekl��$m�DLo�V��Ҿ��링i��;���������E��ShH�����I��c:���Eg!��J5�����Q4������Ŵ͒Җ��S�	�ۉMu�}1<�5&L^l��l"e �(𲲆�	��(�w^��ƅ��N��<�T,��<�q@'�u>E��w齡U���o) N �;�x�e����>Jd��$�X�1^��<&�:��uP��L%z��ه6}.6�k�,�t%w��!)T��Cr��A�q��"������f`��Ӥ���z
9���q?�sqѱq�P����u6��s�u�;�.�nf��?"�0���f�;4ֺ�����&�gK�g���V����K!.�%4�6�ǉ�s����G`}&�E GC�D����fWU�v�$v���9ܻ6�������:�F[��8���jv�E\��>B�8Q��0�<A�0�K,����S�4��Q�l���m���0��h��!��N?�<׌(X�]>^�u��]=���B�7�%����%�$�����p\��f��$�� �m��el�����S1�O�@��48I��Y^�ǯ��Q3��iv�е�CBQ�����q�v�-�U[+�{��G!m�^
5���ض`��X�4�uG���Ѯ\1BÆ:y�b�#�o�,͎o����F��(���)�DYY��+��4�=6�nR��6ǥ4��&S�����2����"<�9��Un���i ���� �y�̀� �y$�1Mr��cс��% ��r5��0�S���~)��P/��dЌ�0�G_�6O}�БЍ����9\��Ż��e���w���^*�i�/���j�(	��ϴ���P��Hpf�(���!B�:P�u���E���O'����	��\3��<���Ll���bR�_FOm-�M3H$�ku3�@��?�T �XS�p!g�W#����Gs
P��0j�w�ĻSIax�g����Q���W���@���c�4����b�t�Q�b�U�T�����]�sY0��5�H5���f%N�/s�$M��ߑ�3��*F7�X�oZ���ɷIɹ5��r.w9)�?qs(���a�
W}P�����2����lBŲ\���j��BOy���c�iѓ���,�����������i->��^�%��j��F�d[=���%�J�-ś1C��M�nn���)������\g���-��G�:�FBdR���
���*%��{�aJ@6s�Zg�@��{���qO��tԛuv*<n,lV����wQ��l_�V�2��jﳮ'�ʀ�/#"ٜ�i��(����U��\��Zn��lx�V�N�"�ch+�qZma�xI�;=O}Q��#d�Zb�9r:�[���:�(A_,j���
;c*Nl����]6������_��tcZ��%��~�7,qx�ʰ�ƶܿ�7�z9���RX���lp��7�R0/X��v�d�Us�A1-@��g�P���"W��[%/��s7M�;Y+r#V �]ul�ְqy�M˨L��B�nlUv�/%cN�a@�r�t��S�MI�a���$����:�u�~����H	�=kﻣ��߀���FS�ſ��4���I����M���:��l��6)w��4�����=�`.%ګ�[�w���Ւ�
R~��Y��WYX��`��/ d�Po��b;�]��y�[~�:����t.	���*�ߗ*�FU�nZ`��+��(w>Q�7F��{M���k�}� �^?YLF��4V�:ve)
�Oo���eoȸ�6c&<�A���PE�C�j)Íh��h��J��~-�rb�-�s5`���}�@a��]D��x,��Z�5��e�.��U�/>�hN�c�Z>�$* �Ii#�XZ��M��<}I�S�����W5�'U�x�I�&T�ۅS�Fϵ(����w=�9>f�a�8��=��c�z�|~݇c=>���ϰ�P��EzИ�<\+��`����v8I��+^t8嚉ֈ̟*�b���A�����o�~G��+�����*�6{&Ҫ.Yzlx�a���AF%~m��;z�0U�ceL/ >��3}X����@'�BzLIZRr���Qlӽ�#��<c��8�\�e1_S��~�,��^E48zE_lݰ�I���Ud�.y��e�-Rj��k(��l�!G�b`O|1ˋ-��$	^��$:`BXJ���{Axۏ�cYğ��z��4d��R���ԦrcXP �F�d幕�-k��N�*�������.�KL�]���U�o!][F������%��2zg�$�`&@-dH���pi����@)\�(�]TrDr�&Y���S(��A	2��5��,��ue���){b�1��}��{���F�����1˿��4ǚ~js"�#7]�P�����P���~�џ��v�e�]���;l��|��\�����:
�(d�vۡяU�Y?�ɾ}h�$�U�gP@᭺�Y�(q�?ԜYS�8�a�^+��:,�`����;���h�JLuT��c�6ypˇٿ9F��m��O��E�����]ͬb�I�w �|o����KܨŖvr�+Y���m�����0���`J���B��ק��4dY���킡+^��]����ɘ��|�����n6��y�D��_^�[9*�OeN�`�LFo
��|��_�Xa������/�H���a�kR#2�/��ԙ�@�0e�Y75ɀ5�9~�͢V.�ڇ&)���1{j�-�,U`3�-�b�88[Wه��8jY�g�R�{�C�_����ښ���@�R2�x˛Gл�����v�r ��$����QmH6&��H��������:��:�����f'�<m|�!��5M:U�o�c7h[a
�����m�B�O���J�~S$w�h���P��yYQm�hV�0)ʅ6��u���!������V�{��WP���([l1{#�{.�0w�)XУ8L���W���D�7��˦��(oq9-gAp�ɚ�҆O��'�-�R\��˾��g2���Y����i��i�D����"S��٥�{DS�Z�5���Q_�D%�!!3eڈ�sG����$c���"zq�=�^�Y��K��.�k���C�G� <j��@� {?���^u1�o��<y�0�@I�a�p�Qt���ih�wĹړ������(�=Q���i�E��ǘ�]��X�K�Re�w2�T��� �����<��=Ih#�C�)J��1a�T�'��.�В���a}HQiG�S/z޵d����L��&~N@���אE���Z�~�͍k+H����ƐHz�'J��x`s��ϹWm�R��1�����0+���].|P��#��~�V$���
R����"���ݛ8�M�g����R��.;����⚘�Bp���g8.h�,��������E�����k=.t8�g��>\����w�燂@s�c�����jG)���\z":�u;����?��)�@)f�0vr�����;��0U�}Z}�e�(:�}��� 6�t��bc��v�?%yɪ%Y�� �iz�1��	�Y��U���,e"�MQ�p-j��y��
=`�E_���zXW���!�m��sf��P�^�@<k�L�LM��KXl�����@���'=� `[��_JzE�]�tM��^��E��#��xX#��+kT�-�FȈS��s�S�c� A`(�9&�z��~[�B<�<��%Ke�ou�۴n��)ƭ��X֝Gy�˦�AdLh�w=��4��)T�1�o+�;�z��T����I��N��^Vv�4$$�2�Hn�^�pV5F�[��T��*�`�#~�.͒'��9�  �[6�X��g�K�� !���'���"�5�2� B7N%cI����X�q�ib��6I����ST&��P^�K�ۘz2g�%1������K.���J<����!���k�Y�UIY����-muVG��!~�H�0�w$y��_�_��I���a(�=�
�䌑����]���H>��e�(|��d���7��:��tʂԁ� K����}4�:�kـ�:��N�����O?g��s���/�r���[�ـ3Ż���b���g��	+5"(皈xW(\R��0�<y�6~�՝M�S!��T�e�����yOM+6�����h��a-�/��}�)x_6�a����b�C��'�8��\zn�\bJ���>M�F�n��7s�O����hJK?H�T�N�0>Y�o}�Y����Θ��u>�U1���.rO%�< ��G�)��#CQ�%G���L'�E����s���I����g����1�?��\��<�g:�{@p�N̆
���'��� �?q��TL�~����y��O�"�dK�����踯FP󈌹�%�q�Iޤ�]^��3<����ZwP|c��ndg:ɵF�}�9l.^�`��/%nb�6�f�X]%u�����q �\q?��a��ƹ	��q~&L6IG�#���\?N�m�jMI�5Z^���?SH��a�Y�`7�Em9���5��7�0*Q��d�����S�	rJŋ��[q9n�ۮ�إA*Ud��`�|zt��\��_L^�j�Þm{@"gO�����S����_h4ZV�TM��C�,�V����� m&y\��Ț�m�CE	�S�yO�T������d����WS�����$�wm�D��� .��}�{���q<�=��  �r���)�Q�ˌNlg$u�H$_Q�ዘ���_�G��¢tP�v���	�7)Z�ƻ��K^\�T&3n��2�D��U�Zl2�v&IZ��֠Z޺�ZaGz��ω`��9mŎ� =BƢ���D/W�� �%���HҺ��A)��)|�䟼�^�w{wV�\X����D�iT9��lE���t/H���ꬪF"OP�������b��G�������҃�l��,�N���=����ru3��?#�"@��W������-�u��V�Yx���'��Ц�N]�;���E����v�K��URo�п��en�-�N/�
�3Z�
���
w��af
��-�t���-���_�7��b��U#�3�ѯ.��`'�J ���9F��*� ^\��<��Iȅ���n��9��d�:��R� 6M�~Ѿ��ۤήz U'��D̪�^r�����$L�Ŀ�+�88�'����}��NR@ܪ�$e�,�Pt�O�T�K��G&�4dHX�@� D �7��U�o�\�C��l�YD$�%����<")��li#*��l��/Q���1��������3]��>E��^5.���Z�f�0�;_�^&z�c��s2���D������'z�F[o��;� ���J}qi*��)�7��ѭoS18}���2LNGO~%�RG�}�_��v�)���Gõ�V��凯��K m�(��.|ܝ��f���Ə<�>�){^=���r$vG�	o�p�*dΉJ3�`o2D4�꠪����3s�����F>M���B�C��.J0�m&'�vs�ڗ�`���s�-�yl��>��y�ؙ��\���ɂ]�����7�M&�����W��M�y�c���Bw�wm������6q��.R�e������P��_V8�M���q&0�
*i�"�i�ܲf�o(i�?1�_Q��p`���K>y��e�F�S" xK�W3��ӓ�����f��t΁W�u.�]�
'�)ҌD�ɠ¿�^��LSLOHr�1Nv	���!t��`��B}V+H�B�O���B�)e���!�*�1��^��C�
���O�P-~�%�!!���,lБVMW�&O�Pn�P�O ���(7�'�_* �s?7�F�v�RYmqj���)#Qa<<��cL���6��k2'a^�h�?���ܛ�#�;z��C����CVs�����	�:�RD�b^�B�o��O�V��Hl;����_2� ��b~,�/A�F����G\�ӟ�"wƈN��hL�Y�ZWW/o��=� �\E4->�-���|u��h���2i�ףR��.�L2�kC?ͤN���o�e��w�ɗɜawmYV���$����NX�yl_�EA���S�����LPsP�g�Q�$M@��}?����܆Dń��R��G�P��!꺐�F�F���;N%<�\���7��#~h��Aٵ��|�NmD-��v���X�}�tɥ����CW�M�B	{xd��c��j��V~��4:�V"(�3�	�L\R]�M{�$�����Y`��(�<���v<�����#հ�x��a%� 4u4��Z�8�.����W�+�J!��E�S>6�k�rz�[v��H����Q\���1Q��x bq�`���,%��8���w�xL��j��s��ya��#�ٞ?��AN����}�8�T�W��WW� �=Q0���}D�����:�n���L��#�Ғ�*-�Q�hw�燎��º*��������D��(E�O��`3�
rW��d�d��ǊI{�+�{�g�/8�r��sV��ز��n�9p�����t\�F�zﶶj���V��<|��K��h��5����ˀ_��m�{B�u��
�c��7 0X�������D�?���[�Z)�T����	
 � �W8K%�q�UãNXe(����%��y����^��&#��t�וRP
��p�Y6�����N@Kx �R�=Q*g@*�G���^^%$XtQ(K�(��5&Y�t[������3Og��HI�xʅ�B�M��\g<Բ��!��	�{>�&�sX�X!p���������b�<���^T,TE�j��Ut�rex9�����v��Π�*@of�:^5�ě������Ci=�N�;�oB���Q-I�TF#y(DV.�ʲ�x[����eG�	����g�fT��I��6p֛�pA�G��p<���9��$��b�#���9���.L�G
�wj��'o7��?����"�y
�)�tN�5֜��^J_��u�Q(�����}�i7�A�U��٤��,��9F�tKҡd�8��NJ��[dPź��9�Qw�W���j4�-������.@�yc��\��:n{i�|$�XlxVHYEB    fa00    1d807F�U:M���6�⮭k`\=���5.I�BC`��.m���JIχ ���HU�~��8X�q�s��u������Ś��9l�w��-|KA��un��55)�&���K��F��4xh��O�F؀tY���^=Mg�č!�N�d�ܢ<L��H�'b-J��r����W�!�>��4�	�?g�%d!��o
G2�z�F�;����	�v���ܡB'-�R��:C���ޯ�F�}p�?o�Z�VA�)ؙ���yg@�ͽ�ap���1��� xqEE�����p��dkd��|vE���n����l����x��8��Լ7p�ܦ�]M�4S���ee{,3��}mR��r��MbNZX� �-����J�}4`���k�s~τ\�Gҍ��ܥ?�|����X��q[^5P �}"�u�'�p�a�x?�KW�A���dg���UH6��Ŗ2� ��%?w�"#�����\�F7�����
�@8Q@rp�*/�
���Z�'����?�r�i�	E-�c��/9&���ܨ1���u�`�7��\CK|���|���Zm��|����a���R�b���ӑ��;	��#�5���ңc*�Y�7�k-i<�U��W� ggh�h����,�`��x`�	���$Q�+��TZ�$ ���ẝ�%TŞ.��".Th@��N$j�4�1�]Ed���g���PC;r�vZ6�����V����P���Q�������G���~�րŖ^��А-:2'�{FX�x�V�c)qT1r�v�l���?Xb*�u[�i�[2�1���DQ>5)��`'���(SH�Y� ��0=42mk�R�����
�x����V�B����]3P�EH`���/���@Fki���W��9-�f�����;*ʧ�q�к�k�Û�IQ#s��S���N�)��r�j�����5��k�YS�\�v�$�8�c3�rP������:1�̞��Z/(h)�)�*�H��KJ�92�ć����;#b[��4G_"5y�w����-����@�3�s	���k�j襯�(y�1����DSn<cM��/��_�Z����Xk�k��I2��W,�������x0 �}�˸��p���x�I["�|�6�3�$�}N?I|�%� ����Y�2�Q��S�j��č������}�F�m�b��7+	)i��е�m�ԛ�L���"����|�a��O�U/��^25������m�
�,���+�ϲ�����p��M���Y1
�:�/�K�k���v�z���^Z�C����{���?�o�lu˲LHR������}g	fN���m��P.�)yZ�Z�Q���Y�wv�Ԏ���d���`I_�V�.1�r�D}�+�jH��>	�^���s	���(?�9�<�������v�e�l�K��X�Կ�ߌ@�MZ	\�a=�̍l�0mT=,����&z {*)T���MN�8�wc�N�C�C��m��׶(���	v�K_E����zߖە��� LK����	O]��N_V�Z(�>jө+!���K�.)��NZ���wޯ�.�]}nf�1IRaB\���͹��Ö|�'䶫��?��� l4KY8Y'����䟝�t���1pqש t�Ѽ��S�k�ظ�����؆2"��H�:Wh��oTs��������a����Ye��˜
��[��Dr�6�fK���K� ��	"��/C#o�Z��b�r�NP�3�\{Q� �	M~L]��fIҊ�D�x�U!��h⃔_��)ӗŜG��^=B���z)� Nӳ7���L�S|,�����	�#��!�0^\jr)���������w2��͓ �A�>{�L˻��S�ӭ�4W�XxdN�s�~ulQ��M,��M�E��j�]�\�BU�@��A��ɘC�T>"=b5���0�j�u��a��i�ch3�qF�A�x�VZǉ���{׎t8�_�W;�W��UEuܝ��u�����O��I�G�q9�.����Lcϕ�ƫ���nݱ��.r�d��b4��ߵ�� R��;�j�J�q�0P7�M�O$ɘPqR��ݙ��Q�\��M���r������-�����}.�}ÆA�I�I�\�w:\P�C c�ԕA�O�k'��& H�sV���x�Dm���"��?*��!�@,�2?�X����B�VP�̚�=25|��H���2� ���n���R���ΰPn�����IewK�U�拾(�)A��W���-��ThG�������l� �'2�it��I����fV�R�	��x��.>�.L��6��XQ ����c��˃�n�㧼c�YQ"Б�c�-�+�����q�+[n�x��V�-�[�aD���+=ݚ�j�i����	(uz��}D`F�a7�L�QW��,�h��,UԲ&#�GG��)9���~bǱ ��8!\�z�ՏM�\X�ྀ�)wkhg��%ATO�sMUr�*��-q��̕�9B�z�1^PFy��Q�\�K����\bc#����Y9_���}�Q.P�'�B?gü���� �G��%��F�@��n4W㛹:�y�`f��9!�e~b:]AF��o�$u1xYs�J��	�T�G��Z�j�D|L��;^�Ţ�ݞ֣1���OE�tI�6�α�/��ܭ�t����}�]4!��曲��r�̈́�+�D	 �e��;�Ŋ�; kM�qaD�O<Q���{٧;�7�岄tt�ۨr�:�}e��!�;�S5�0$�p�~]��7��	�$�Ue��Pِ"Հ�g����$#��cX�$h�����mʿM.5*�i�ڒ1���"J���s�N������.|}�)J2���N�vl(?���|�$#��,�3 R�벨����g�Bg�m�d�Җjz�܇k�槧��K!QW-��R8��<��*�K"�A�'��5�N!�A��L��!� ��H�6v�vDW�`0^�=���a�{�,��TH�1jןs.'�K���l¯3MQw�M�WH 6���
 ���` �_}�,���R�K�3ňP��V�y���iҟ��u����lX�v�"$��|�+�c����F*�,�ur4r��&�ĵ	��qM���&���I�3��!�-v�.\#������lSM���r��.��� 9��<���Is��˘��7����M�&O�����6:ؿ9:�ld�u�e��\G��4[��XԪ��tC@��c]��dG� Y7�(�ø u�����uz2
@#t�]y���^�k�}�� �m����,A��Pf�I�l+<�p�i���n� 6FΪ��� �����JxF�����p2��B�sد7�T]`�p-�;4�y�
�Q�}�?��&��dJ*Gɽ��{N�^��W��衢Q�IC���Q}9N��2��}k[x��������m��є�UL�3�'�~=|���ե�M��K�p��P��ZC�e^)����"a�2P�ŏ㮏wݴ�|L'�W��*q�ˏ^>��� �����	68|B�L��Y.�:o�l�l�s��Yo�]�v�>Ƅ�37wA3tW@������W�]�i����)�k�$[�h^}/ml/���"����\�b�zB(���۴$�Ǹe?��;0fكo���x�����v7��F��Pĭ]_F�Xc�\��Y�����G6	
�	g8s��������Kn��sPؕ�:���0���K�LU$X���T1t�)#dt��+E6�?<�f�)%��Lk�oS.�^TA�bg�ݹ3�ޣ�b��9N����8�Ì�s<�͛x�]���X(�����(O���pfV���s#f�&^�����	1۠ �����a���_��sAҺ�S���'?�@�֬���2e|�X�ѫLe����d+w�\]s���6y{�����[��Tf�$W�F�y��QFl"��ܑ2�tN�	Rق���~�y��̓��*F�����h�����]{�
M�S�#��8��-�F�@1gC v�@&_�ql)'2���,O���%�nnV�(Ǐ��|#��ڝ"Z�rTfy���׬@��r5˟)�~A���̀UxJ� ϭUG�H��Sn[��ا�@=e���,�*4_�;��6��;iJ3%���<��#o�'��%��2�:B[B�oM;��G�����g/��?�7�!0V�o��>@�:��i ���9`(U: ��Rn��
�ݪ���Xa�.�,����:�0!)5��u�����ʹIH���s}���yb�Wl:�!�����T�>��0Y�a�����wB����ФŘ���^�4Ẇ0�(/6!�(����BYe. �'�ݤ�oB���w�o3�_x�q�^�ˣ��׾�$��u�m�V$�S�\cd^�)�vl�"��F:��6������:�4g�B�`r>N�>�.��Xa�\�gzTPS�W������%�\���K'j�u�EP2_�94�)ʥ%+$�X*�����B��]m���S�yG�yh�{���al媝zU
G.`V��	�
j��T����s'�& (��SD2�`鍡����E�Loo���,�����0ٵ/��Z�_J�H^��S��1]�R��oݦ:W�����2�n�f�2�l��;��ڐN+E��le5ت��.Z�}7�(G��~��>+,�n�N,/I���ת�4�.� ^ʾ{���Ac�|^����7��[���x�`�P������̪Gݚ�x�T�\W�� *��V�g�[��,R ���q7"aw�IoX�߃73-��2*'��r2U3���J;?�\.N�Y��"[2EV�{\��O�Ƶ�W1���,�J�؉�?j���U��}v��L��{=^hƐ�[˷��\��j���D�)��i%��Rg�:Ʈ�r���9`L�p���S�%��]a���<ݪ����~����z�y�}��j� 5͇��]����f2z����4��� wS7?/`qf�R��[HcN�
�y%$��o�����:&��^S1�$S��z���.2�bGi�ɤ�`ֵȑ3q8��'�|�xV㐀�q:��i5��&TA�f56 e�*�~^,�ۈ)�βRkO�\������uA����
e�uz����H|�����ny4�7BI�*?@���Rx\]� g�	���Z`�S=��üe��8�H=�j��GK�=��/}�Hv���腖�G�)k��={߸8���T��ͫ\
��'�'�2�0#^���܃-$�1sXaC[�����p;�u�����-N���?`�l�[ �@M	.8����5/�:�
�Cj�۽�s��JP^���%�u�!��un/ ��7�d ����=��Y����GWR��x`�����M��:�����%�����N>��-����V=M��5\r�$��U4�����,�\Š��ϗZ�)Lɑln��TE�m@2�_Y/A���r��k0���i(9O.�� 0�w�M��уSLf��%U��*���{M�l�;�A�%���vs6����_؋��B�K�r&����u*cB��Z�'�Z��2��X��cx��Y"V���iI��Ϯ��eT*1r`Y��������" U�5�-Y�k�uU"}{e!�(�j4J��V�ps0�%�S�9�G�~�uE��0�����*+��3���J��C|��pΑ9����p2һ���@g��|qq���iM9%�n��h��R�$ݷ���x��FN�3r�`r�2	�TQA�2KYF��rՄ�~�h,fT��Nco�2-�#��a5�)G��J���)�Z�+CC�-1��i������'5� ����ϵuW}t�ԅ��uCn�C��?j�>�7�D&W�����M�}�z�v*�H8�cӘA�?̭?�e�%�����{d���n��:6ڂ>Ehu�3���q�$}�V�E������Ej�6lq�+G#[�W��%��K}�W�y:@�7x�<�Yg�'��Ƅ�$�S��M��͇�m�GNR���B}���'�>AUl�~W��6Z_2��E�bfo�a�k;��$�~��o�%w:�����,��
�9�CRɊ3ra5T��A�+�Ƨe{=����K���3/|ì�0�а�k ^|�X-T���%��h:��;���������xz���K3s�pǙ�q�˲�rIX��㖱�h��]�Z
i�j
��K�ݢ�;J�m̐���	�f��r0!a�I��õ��y \
�V���:�)�|.Hy�g^9�i�~�t�,���6cq��Y%�5ЫA�h,�2�`����+�C���m�{�-XG�H%�Z�o���R�@�D�e~��Ϙm]�F�7������[ڛA��1���:
)z*P}��D�XO�MB ����r`�P�1;G��q���3o�K$V���m��k(њ��N�u���cq�)�~������[�jp��,xɨe:�5<������eR��� �s�Q�-�&P]��(�~c�����E�p�pZ��=��<ݒqЅ�Ԫ�������4�ֈTNi�$��n5v
�����6�.t:�q��/؝%�ǑAf5�{�J�tO�S?����Y�PS�&��A.�8D��*p'�'T��/�r)*�
��k�W��ƾB[�TM�H9;�oS��͠�d��6�^��f4�ꃾ��z���pT�O�A��5�k�|��vx����}����d,��g��y'�j��r|5���3m� �q��s`��[+R����C�W@���R���|�!��)����򰺤�-{J�t�ǿ. w!h$'f�DI���fm�ϧ�p����p����g)��� ��Tg���z�{�0�-���Rj�Ymɢ�iW�J�h�C���!0�5?��KW�@�CU^�{q�_o���!�u>%7�u'����%gk����*��xj5���v��zay� ��@z����'�7�R�%H�o�4��#�WWY�|�p��O��m�J��R)df�$]I�8�!+&�K�Б�J�c/=�V��/�Ej��$�O�O�`�z�1��$]�M����"R�:��3ż�NOD��e�mT	E�p�F��ST������PbVipN܄��3vFV�
��*j�v�:/��L&k����@�I��v��e���C�OKP�9��b?��/+/��)5�k�y�Zc{��4<�i`�05`���ޗ�O+��~Ġ}K;H���
[��r���3�]�N�~��K{�@��e>Y�'�<�����	�(��nX�$��Qy'ظNb��<�=��#T!<�wk�2�ƚMH���1�f�i~
���`���`r̛��$��V:`����$�����̫������7�!����� �� �>�v�6�]�'�ո3;�l8�1�y����n�R�<�}���	����bG}˞e�9<���rv�L(��||���PZ#�.��z���K�����XlxVHYEB    fa00    1dd0~�u��C.u~��N1v�'��S-^���p��l��u�|2��M46CF_#�2b�$)�E]y��[���1q�?����O����J�F��\v2�T��N�H�t���Pٗ���,�x��#V4R�!9^_E2|]�&č�,�q��L����d������r�?g�j`��4�F�>��\X^q����]��2���~EJ�U#<�Tw&���o3���׀�<�dZ��	�62n�Z����!��|���Q����h{ 2��	i�.��p)�V���1�?3�sB�lf�\��P��3��y�^�a�����ߑ�o�Cazڨ]a�K�����Z-�k�����K��!�aҎ�$@@,���.�K9O��29N=��m�n��i#�n���Q�4{�[���J�"e����}�Z����ݡ�@�ܤx�*��N[K��{郠��.D�N���ˇz�Q�zýa���ҷشci����S�/ �㯌��!���j۠j4�by�;����w
r�M�����,��vF���kO�!�����l�� 0��+�{�UA�������j�����V�RT]6E�CS|���=a�GD��l#@w��W���9���&_o-��G��3�]���dLo���|�`�F1
Q���4�͊��t���DGPc"ndᄋY�9^�T��^����S��m���Ϋ,a���пGʟ�GZ�swE�~a>���	}^1�6�N�"�+�D��I6�q-f_���}iE��&�]0~�X�Xa�O[�W��#{`mVDs�̳�&_��ۉ�TүJ�2�-�G�����Ok	�>Lq�ʹ)8>Ӹ�>Iu�+8��C>mg�2w\��������dM���X������/�n`K1���7ƺ��/� P+����z�4�N��FatB#�ư��o-�"�Ѩ�w$o�Å���ۨ_xٱ������y��HMю�r(�V(Ԧ��Pw	xY���.���x�Ncw}���(ęQ��Ze��n/��Ghy�bԇWW�Z(��Z+����������iMf���H�GF�1�X8���$��R��|����y�4fQTt 1�Vn�-�&w/˟P ����.��}J�"Էf�,:Xs�w��������f�I�"pG��<���4c	���<��lf�U��Z��.���e�YZ W�T,w�Rٵ* �*[`����,m{jq�b�("[�>7�������`2F��	U��)1-fK[�c�/��s's�)�Ǭս��ZU>sf�rh!��Ӧ=o?���\��� ��o�\SL�~M[F~4��}E|ϊZ=dr
����b�@Ϛ��u��O���A	z�9G�.��fl�����/:+i{��<�iO+A<ַ��=r���.;�����;�E��{���L��:Le�
tײ����Yf0���^!*������p�Z��!inu���
��y`����_�:L�5�0rܓ����ue�U�@�i�2������Ƥiu�Qޛ�(�HҒ��,��P{�D�u!vuNr��) ngR)��U�Y.*x�("���`�/�̌�7���A��9��D��qV)�����|+��ځ�]ך����0i*�l�9*��0��'���!��>���'.�q|jP(�5��;,J�<S.�0Q��H�_��E o������k{�'�v�M 3Ҍ_Ծ�D5���Y�/]JIn4R���/�b��i�4�W_�Ё��#���Z��N����fQ▨s�V'@����>Cd�d5�tU��R� \5�~�M�vX��e���}�����ѐ��I
�(�B@��Sr7�&�됱�𘦑�'�C�z+�V�]�H��D��׍�R��Kf����.���Ha���&���3/�h�c��Í�4ǥ��4J
�xz�l;�X����~i� �6�GAh��,YL���A�g*ê�3�)Ĩg���d7� ��Q�9djNI����&#�՜y��{�"�f����@tv8��8%>4ҁ犧C?o�������.�?��y n������{i�*����T��ugi��1 ���eJ-�{7�f���MJ2��:�9��'�rշ&x������8���ǁ?�Z�kbLFLp�ǿ��?j�Ыa�gM-��o^~\U���6���'�����~�l�wg)�7 Q|�|�S�ڴB�%U���!@����o0C3�0�R:r(�P����Z�?�j�H]O&��<෥���o��\ڠMgr"��>.
 l4���æJy-ZpS�?���ac�h�o�a5gU���?�]�A?a���\l�T3��6��mV���L%"�k�,Q�/־�{8K���v_�Wہ鄻�3�o���, �ׄ�5�2����'{ ���m"tW��ŉ������0���v�j���%ˑ��!��~j6X���?*
� g6���Ign̛+-�֘XI�c��%d��v���q��k�:��*Ow��n��0��c4�<<X�3G	,����y�w4�jYw9K[̘�����[c7��c����aj��ĸ��ˢ'�;���7k�g�`�x���ό�����T5Ę����� F�����.;UG��#��(I��x~���V�PG`� L��*���Z`��ݺ���\Ԭ��B� ��b"h_��|a�\<t��;V�mn>Q�v}�H�
�Tu�,��kĴ��Ю�v��!�q�|�^�2+��ɭ8|�$Xz>�r����	�Q��ZŹ���<�%�7l����*#��g���Y��%��`7�mxE���_!�ݾI.�v<�eo+T����q�bό����H��{�
�2[�Q�6�����G����ے�TÜܓP�B���j�����;�|i�;��=J�gK늊s������{e�~E�&����7�0���H����I
B'��Z=���O���Gӆd��ĶmGX��A0ޮ3�/*�9����a|�A����/��å�tm,�G2���c*�'k����L'"+r0���B.�� ���
6|�t]����۵L�
�,�R�Q��ׯYw�n���1,a��&��:�Wg�)2����=�[�y�7�9��c�抱�4A���P��y�����6�\q�6�%Sx�J�x=}�M�L,���.5G�I�?	�K�8�(�m���ܰy(k��a�I�9�<m���*d�A}�p�ׅC��?�\�i�D6�k��+�ԽK��!'SqY�&g=r��ޢ��֎���Cq�A�܊�Z<T9�է?��r:�$�����V��aܙ���n��yC��3bE}�Q��U��&��{�2t58lsi������J�W��5S��"�j�����wN��n���ൾ3�����RCp���C�b�T��Գ��r��sw����4MM���X�?j�����mbeh]6���ɍ\4 ��Φ�3g�3�E���	��V,�b@u��7��� J�;��9S��`@T����$m�KGЭ�)���Dmye�
&�A�@�d7w�8���,I]�,�G����W��%Yݝj46�2�������Nܰ|���8!���'�rp'��~���X��b��)���gD)0(�1j�<z2欀�Y�.k��i=#ý��6E���>��è~<����/�=9i���ogEvZ�?,��^�4��x+�4`(�YM��UY�ç�eG���VHi��fEsx�KՀ�Zv|��3ă4�Z �FR����Ͳ-ڎ}5�y�ߴ�����Y<��*m���+�J����-*N$RzY�����D�x�`O�d�w�o�����s������%�d��Rm�fV�_����+O׹V�bd�w�ɉ�'/+�������է��5J׻F���Z��~<�D�x��1Ѵ�@�ͤ-���T����j'�(K��|l
��yX/��h󹌢s�2?|&-���k!�ϕ��+��=-��q���� ����ŷ�������������ηw���l^	-�>�CгD��(c����zP�u�-��C�:�`'�T� ����rt�t�Ҵ_8�{,^��1a#/���J������r�6岖6�P����r*YP%�M@~�ey���b������~r�){�P�U����d0:�!��;��.��h��w���~4�*�SI?x]S��T̬U
����<���?��h���c"�uվ�P���xe��Y5,ݙx�& �J33`�i����(��k�W���s�#��4F=��ԫr��{EG�x���d�+��H#��<�_#��{$�qNI�N��H���؈9�G�wG;���8��B|P��w�!F9몊��|�0]X"=�SR���a��q��{*(>r-n%��|�PDu X�^,�?�Q�f��R%$��61좞�ԍ�ɞ�9��Y����m�����Y5t�.��Z������~^g�W�Ƃ�*��e����ҩ���|��)-�D&�e���#��u�|lzt�"��Ax1�ɽ���b�-V}�O7����0ت�E.�hP�N#/�]Vh�S�/��訩�|�$5���zlr	߳�$�qF\�����T� 5wed�@��ӪM��-f���w��(�:�~'��y�'���5L��Py��d���5��Y�qw�?��=I
�!G����ۇgڋ��S�_�-K�?*�w)��6h����.L���K���ŽD��Y��aj}�F0�G�dx��b�F�ZPy/xIҳ�ɍ���;�{�~ޙP��mz�	���8Z��'5(nx}�E� ��,�~J1��U쪝&��"Ņ�������uS��2�@w+.����ӥe	X������"����g���U��óbZ�ËG߾����!{u5꤇��ol:��L=N�����9��p"�2��s�/K����������Qɤ��������J7f�)����d�����
Jp�a��(G��4C��rB�/�sL��S���q�����C�Uhd�pr�O���E���f����J5�����_�t�T�5���XI���pW`�����*��c���������l�I�Cx��Acb��p�����B��7Q�~i#2 fէ��7�mчi-͖��sD=I�z��;s �B0Ä�rwM`�c�K�Ht���S��ߪ,���\�)�Ɩr�Ͼ�']��Sq��l��E�"OY^�֚�8������Hw-�/�8���;�nk������u�z�=�F�g���˰��|B8F���(2����]�?��>��D[v/�����X	bC�Fg�����3��Ғ�Gv$�Ե�`#��}볦͍vP�aڤ��i!�������B�8�^a�?-b!� ��a$j��  1r��1��9%}O¥��R���Ѹs�A���B�ch�03U|�������e�K�`���%�Z�" J�h7�<����uA���'d������/���G�$b����T�s�+*�6>�ĆE��$��&;�����Vc��@VKC�T���Z�tժ�f,ɻǿ��W�`��d{���%?u����.��)��� �2��)���d������p.��1���5���MO����V��k�φ2صti�˓+b��wۃG��Z��p�0�zS�I�W.<�C�W�}"}���y֣,�c�e�0m�1*sμ�a�Qb�eLS^�MI$�J�c�l Ӷ�qiʱB�1_�5��F��0����X����UGʐj�i�|�G���t�J��3g�:����O��5�!/�/��ơ���F�~d��L;���$;1�q��Iq-�΀3��έ�TBR����}�~t��ݿ����+�8���qɋs{o�Ւ�����6�䜠ƀ.�-]v��{bZ�lVK��PT��;"+��=0I��w
�>J�@W�Zâ@V�_�����P2:�u$+�����d;Om� 8T
N�Hj�XZ?���Z7��'6??!�)���]ŕ���M�����Ϋ�5B\��+3��C؄"C��T�"��U����Ij_�7���3bAH�΄�-�+-j7=���#Z�ysj���/���tbq ��m�߫F��p	e�~ qYc[���Ϗ��Ӷ��,�.t�.9�KŊ�o�]�f, �����"�G2{�\�D���W�Ƒ�ш�ߺ03(�3���i+�[���nruc��D|x�B��:�ν?�\��нA�R���O%%��a��5kutE�W<�kA'��y�j� �'̢2z*%� 7$O���y</PKT�3�,�:��rT�YC�;��c��e�X
������ֹТ�xN�קK������se��_6ETt���VE���]ǋ�D����H,��=�Dk����0m�bO�����o'C�w*���b���TgJ�(zN	�s������ݪ��L�~�����|�b�K���YO摘�W+�1��C���:(~�SPN��cPk��
A�|��5kT)znEi(r���NIhD�д/дm9ئ_�2"�r��^4TB��*�&�H |��#���x�=�/4�J���L���W8�r3c��z��^����h�c���Xh�#5>>��}x�D�2�6|�-mvi��;��=��#���'?K�$$��Q`m�H	�@�/���Ns0%�k7�b��%b������s�L��m�����+�� �5�\�[e��gh6�WW��߰v�n�|"�W�c&����"om���<��̵�&
f��wa<3ȥ�����*�&f��+ʯ}
J�"�'V��{�����<�L��;�
l���m�H�@�|��u�p�\�Boi���J <�+�U�RW�_G���[?��16�6m=�?�J	�����Z� �;�Q�h��J�$�\��r�b���f���Aн�h3�1 �0�� _���
��C� �'�Vp�Ihl�ݏu�y"����[�ۯ�3��;J��l����,БY��+�4H�S��՞�����9͇Oav{�v�Sy�z�v#�U�]�YI)�p�ѕ 2�U�m{�*�|�<��FxP	�_p����Cj�i��3�۶�}�j�?�a���Îg宏^��|�M-��� 8�%�_�^�G �Q�g�Q��V�}��hm��?�ܗ�''zAm�s�jH��Ⴔ-�.�:�_s-�ǩ�Eż0�]�J�"^a�'�h���Mt������:H�����{��]rx��c7zw!>@_�V�S �^V�a�)�Uz�9�vJP����1Nt���M�����AJ���8��ϳ0���@���q�@"��R�e��]\̛Q�G��6-���S��F��d��ZP�EŜ��]!�y�eu|���Xc����yٯ��oz�Eq.]����z2�*�Q���w#��y0+Y�����|wD�TGL�\��FV�����m��!`��ՑC=��3� ��zM�("�آ��v�`���|0e�F�}��)D��|�ό�����Z����3'B�N?Ce�mg۹ɫN���H�6��5~��Gm�61XlxVHYEB    a74c    1290��E��E�f-N�s����x����K�T}�1�ci= �N9t�1xZ�rV��`8 l��-&����f��m#�1q��)�q:=�$J���tKO�z6� �~�����9�:}��O�Jц؆m�qO�9cV{y��
���>�i婢�ӷ�����S�'�t�(�l��|�/�	"	Щ�1<���c���뼜9��ېWP��3Ab��J!������U�y��X�?�n���C���/^
�jU��c�D�$� ^���j��N�����~%G��4�u\>�ϚlM!*A�AbiT�).6�k5q�[�6N����Kڬ�L��o�E�4��5;[�*�E:=��xT�q��W�5�_�o1�&�g(I�W>�Z��Y0�B��PB��i�U��ݏ+�;�>��|�� �8>n�J��$��:W�]�z��ݾ��_��R�#͒�P�")F�F?�ٿ�tV��{��A� �Nӛ�Ơ/կ��!l�,~g�K�T����BE1�q�x���!�TN���.
�`CՀR���sw�������y�M� �Oꪳ���hN1�h�	<���]�?����?k�����Eg�pG\ԗ��Z/��6��%��6�\���
ߒ�p	6p�S�a��Q	S,�4B\���!��E�
�a��������!yJt0�ы�{�m��6�֓]U��W���lC���]�,J��
����W����pȬ��o�V��*Ñ
�W�y"��� �iȬ�v��7��eN�����*�D�w�Tc4���x?����}�ɞ$uw�3�:�l �qƠx�Ĉ�����%<��s�9�p���>��?q�_�gg�$����oZEx��k�{�	��@)c�Y�E~�Û�V���6{�N���"Pa[�ى����Y
���d�l�?��3B�~oA�N,���K,̗W_R7�͏�F߳�I���]�n�W�J���ζ�5��-��R���f�C�Du4�D��g�=��ai�(C䬉�# ;Xq�C��*�D����X��K�bd���|�nHE�_���!�l�RB#?����btlhp�bZկ�*FUj?��,�"͌+���J�_���ڇ?V�٦
�Z&e�P��eϭ�����r�	�-6;�d�{���b]E�H߮%C�I_#e�����-�yN�ڗ���\�G��kc�k`�R�:I�=˽���:y'�w��N�9����G�Hh���|�?g��C����up��N���.���ǲ�ݨ�A������I�m��Y0$��&<-�Q��̏�$�ߜ=�65��:@ �t��g�| ��H)Ȗ (���Z.A��벁"����_�$S�f�SA�Q�(�B�X-�Ҁ�5
�("���#�\E稼/�R�����'\�!�OG���f^����͉��(3���5R5����0���;��S$��t�~��T�^B��~�tϢm>?���B��ך�جU3�(|5��]1�(�a2�\��	�k��߾zB�O!܆TVx�D=&ý6���L�'#���P�C���o���mp����uk,��M�e�n�򼉙�([�2a�/v~n�~Y��0�9�d�{$�	���!2�%1��C#C�*��`�DWǸ�>f��oG�_�`������]0�ML3��_�e���9� �:�`�c�Bw����v<Mq8QS{�o$-�[�t���K�E�1����{�Nd*)LU���h�W�m�(3�>+=��1�:�4Ъ�_1ӿ>@6��}��^�ͅFO�JN6�5m7�S��U��!�\�<���p�&Sؒ�D*��E(i� ~�ȝ\�o�\�r�.~]����?S
R>��׾�lpO��*xۯ8}������Q���6�6���D&�������z���C$_���+�,T8pT��_0�o!��5]�Z}|�c�(OD�&b��Z�`ϜŐE��&`�ho������&l/�B|���Ȟ��~�TL:77O�7���w~�e�(W�i.D�>�1�D Ѹ����oGV>����,O�r�(�Wz7��ss^��֖PoM�������6�� �q��"u�B����b�����|�૰�g�TtEV�9�qK�%6�~o�Sq8l9-0�,A9�Du�hu�t������ȝgP0/���.h�y�T���Gvg]e�Y�+��5�  i��D��6:_р{%BG��/.��nN���	��`�{�P	D�䷫�]�%l���c�f�AWSc�h�*�;�ܥЊ	�dt���M��XfEr�!.� ���7��eE�P��� �����V��~}q��V9���Si���mӻ����ˢ5��⋏|���󪣇�� ����,�I�-֒gǎ,�4���g��n�)�_���ҫRp����6g�O'p�����3�̥��%���V<^`	����}M�`ܜN;B�hp�8~����;�Ȥrjz����c
�Рo��:�,��d̗H6te�K_=�c�6΍??-3��.���!X����xw1�$q��N�y=��V�w�Q�,�x�O�&���o�& �8ڑq�X��K	��Z�
>��nޟX;z�[�>���\P��_	[�ieg������H��Ų-`��e1�4�P����>��|mɭ\�g��n��ba���F�(*z�IְxL��6�-Q@K-��)��]�	�O��.{H`���>D���|��"7퍊)~r,������u,l����Cv���Vu�v0�,�}:%�w��."�=�,,����gK~����4�SPo�vW��n�i�iU�h�A�� �R�����'�����D�6D�C�:���G?$� �ǖ�>�✂��
b�g��pAiXx��<`]�i�n5�Q�����B��� ��jS�/����3��*Q���!eio��a��Y 	���ə~��w�����L{Č+����@�İp�5����m��8q9��|�A׏I��Sؐ�N�K~��n���y)��ԇ8�L ��yr,1H��8t�Or��ul�%m�^�D|=�⵶0���7G�2�,�,�T��QX|�1N/����~��y����M�S�rK���WC�[�
vY�ِ��
+�=U⡋�)4Gy,g`�-�����仰��O�V{����)���͐9Ea��F�JB�<��~�B�%�$#1�qh�"��	A5!�H�m�h���'�����L�Y�C�j���<ߪ�#��1ǒ�����B}n�-��Hg�CL�ԥB��NC�h���<œ%�&r�=�b��]<0�L.���/�A'�}�۔v��\l+�A��Z�C��Q��P���o#�NS|�5k)���v�T�2���y,t�{��[�;%�s�-훐^�hN��I�,G�sM�c���0�{����zVImژ�٫�����-ͷ`�/̔}Lzg��E��6�8��f6B6t���IIV.�]��#�	�[��K32��A�I1DA�RtDvڊ�Hk�&�-Dy=*����&W	�*5���| �b����&XKգE �}�G���zh��l�QuL��1w&��'�'��*��`�ή��\}��uf��OZ9 8���t�w��^5�)K�o�W8��ua�Jp���A�������"Bo�$!�9!��/���]�U^����zs���Uft���,���J�8t��l���f	'Ix��PЧJ����-�
#\�@f����=i�VN	:�b�j��=Wa$�9�����S;��g����r��Њ�r�έ��n.��J7аN��F"$����$�SF�H$	���.r'%q��RE�K��h�K��a�:�N϶�m%�v�x�9�_�p�t��}����ͫPSOz���i[g׋C��j�'s�ɡ@8�w ����4��7�� �A�y�d�=�O�6\y�%�렕΃n��'����Q\o,.$Wʥ��n	�౸G�z�/`�P�W ���*(�����Bq�ʮ�����?#B|��Ia���b��qռ��^3/&) �C��¡y�: Ac+�a �M�b\�s��G�.���C^�W�,�-<�|�C�#�5�v��`����쇫�����&�y��IÃ���H �DPg����Q%�[���C/���TV���PMH@@��˂5�~Y3��ei4/bB?��DI�q=E�8F��F��u�z�5M8��<��kS5��ҭ��!F�W�Gf|�؍<���*ae�����HS����l�=�8+7@���wo �$.�<#�����h�����E��u�n���VB�OC�.e����l���4-�S��(;@��2e/%��!��(��6�nr� ��#D���ҕ��٥��dE6VE�߸�^�S��G2R�w�E�pv��zb�Hr���l�~���7R3X�QJ���K�〨ݟ��9c�D���ξU ��~�n ��s]ݚ+���tB�b����)����,�fTJ��v�,q�bh�O;VW��\��꠺"T_���n���̯�|! x�û���d�8�*ŻA����ߎN5�׫' �ު��+c�e��$p��<��oK��F�I4y���v�?6k����B��H�.]2�Dw�X��r���q�����"�J�M��t� �@�G�����G��9�v��A�ép���q�G*�FĀ�'6F?�6�eQ{a{}D~o��