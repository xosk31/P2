XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��w��i��	�����C�1���wX�J��-g-.SH;��Y����|�� ��l���<��:O����V���"ϥ,�7~��{����i�%�(;gq����C�^5@w{�\��S��<˛&܊CvE�mfk ���\4�q��r��h
��*�+%X*u��C�$�NDo�EV��
`'�r��gFN�"�r46�h�ws\9��\�{`���/�賔b��L����'t-�g�#*~�~��d$��.M�C�QaX�)�|ǧj��6S�[�4�a�+\H��E�xbf�E��W@9�����GŰZ
Snq<#/+x�)��m�Z9,;����υ�t��n�j.@�����$�nxK&��aV�k����a�#�������g��x"H�Y��ت��ӗk5����7�L�K2C�_��\�l}f,��|�ai@�XDl=�-�a�+����<�Y�S�A�<-��z傒�2�OpʽWgƮG?v�p,�wu�ނEH]��\'nr�o��ss��8���_/<�,6G���q^m �>D��2׬�»�J�>��sk���]|���R�gzr�����!!}b�g1$��aL��p��	��QP�란=�dX���:Gv?f���0�.�e�$��c�?��W��2��k��H�L����nѮ��K�+�Ѕ�O	�5A=P�@�KB�-�_)2(ˌ���o��Y�X��W3���2��E��<��%[�E�~ۮ��3��2� �)XlxVHYEB    2bb9     ad0�O���ft�/��ǴĪ�� L���=�ΜS ���� �n��#�"����5�����
a�;ke�û.G���=�e����(�l���9N��I�B�,L�w��U��ԑ-�2������\�| ���e�C�Pv�X���4�����g1���4��@ECX�����'cP��Д�r4�D%@����}�lcLۜm�Ar�lT	1��m��d�{v�1s����H���;�(4/f����J3)$	�x�/��o��pcNh��(	fdY�0��\�)��!�_Ǒ� ��r+�b����f_b;�j
�dMSz{咊�6P���iK���)�~�a:!�@�N�bZ�A7F$���3�A�h�I)��V,�����I�}m�����,�� <��r���S����:EUdUj����ĕ.���zj�b
��(��x��7�
����y���c=9 �;�|��J�Jqj�al�FO��=�2�Җ)�4��@�gj1WH��a��L>�SF��#�H�SǼR�U�ԉMە�imf�P@?:���A�Y�����:�3B��?�U��Hz��j�W����L��{E�'��&yN��@���@۸tw��zo��î�0S��8��+�[T�9�.-��iQv��/�%����o�m�l��6�~&�}���Pj��;�#�* �u�@@`�椁��,{�P�Z�X�&���M�9�����~7rlGg��K5�.V��N����߶��Z��E����q���Y�8�b�n�&��fF`�/��E���V8�|���3��Gb�	/�ԙmO�5|���K ��X�z����#F!}�	�EO�Gx��+�H/ު��>i���r|���;�-+<�G�,��v�H�sn��"������t6#9�e?�ſO�T*�J63�S>`�'�j��(���$$[�^z�i��5:��ˊ�v�qFI!��Se��#M���y*��WUǋ� ����}j��z�,��S��!
�bR�8�A�hHr蒞/_s�$+��L$P�Ѵ�nq ��G�Y;c���܏���J�6
:H����\����-2�r�v砷.2�}-�1�y����y]jz��X��5 ��&���Qn��V���f���|�4��Y��jZ!�#э������ʺ|e�Q��Ƕ
.[�ۿњI{�A��YH3#��B����b��d8e��&e%�����4��(�L�ƍ���g�&��w��/�(gTK�:���8A%�����7է���$
�Ioؙ �E��uFE��k���8H�!�?XojR�~b	ш�Y^�0�vX1~�J�|�SplN4mq��-FGō�}��'Э��8�j��lE��1����x&�q�MF��^s�ȷ3���0H"L���@/q���N	�gr�V��SP�Kҽ�$F9�(�m��Wy�D�'�H��D�� &�}?���rT��͢+Y�1��T����,�̈B�d1W86��ٝ����8��:V����>j}��}an|A�7���"�]�;�Y�(P#9$�t�F��(ڰ��[��:�����˚�@��<[�c�l�e�@�n���x���� '�mR>ope��s����G��7��5'���/��HkQ|���؍��{�E�Sb�S�-임ie]�iQ����M�9E��E�@��0��1��_���}�y~"p}����zoч-ʞ@3��yRE�Ads�XRΘ(X�G� OO�s�n���W ��7RD�6�ތsژ~�`�(���[m0����HX	B�/�*Bz��;%�C;�K�����$Dvs�/����p���״QG�ܿ,{�B�H��hx�>������b��x�[2\��0�ޓt6R�����IjP=�mbc[M�&����xFih��h��j �53=�����o��)��B^f��|=]����B�����$x�h�7�q�S�f�G�L�_��g��#��?�άNy��0�K�!.�=9�R}��[AIhG�����'�X���o5"���Y
�_��ѓ�Wy�$�����%Kt�5�,�A�V�4��5�*�Kȸ��LV�����؆�όYA�l��&3����ST�A�e����,.�����0>�������/�X`~���Ń{h�f'_"ߏ�QEΨo��y�����6�����~�޹ ��۫��|�d�[U�v��ܸY�w�9s�Sه�'̷G�G[�`�������E�&�[�������/W���r�wȿ�,x�w�4�qN��ۀ�{hs�"�oʻ��_ �#!,��ʛL_�JS
zx�(y����e�~�먁x}���>-��d����G��+hw�+4�,��v;;B��\g�t��=ϕk���_`~Y�+�����I2�E-��h��n�
�M�z&)Y�j����#w�vL������%���V����:���,O����|[c���Y�Ք�|>��$�A�k��k�PBA
fQ=S�Ԝ�#�|�;DZO������CT�p��s
`�_����K�l����x`�|���P	�I�w�z�/,dZ�Q8}�7���nu+vC�(.�?�@�D�Y��^T�&�˄���z�A_�:�q\ҫ�t��Sr�r��'�m�U��y���.�*�(,UG���)P{�dSvA�ȿ�씙D��������Ū�	����XX3�Lȿ��p����v(��[`Ԫ2�KD��a�п�G��Rd�,�*��GI�