XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Rt5
�f�,���L뫿R��?\�h�l3DjL�	�����b�b��U�l�;�TX�A,Y��p��S{�=�#S�<7���v��+�2�Y��Z�iJ6���ᘪ/���e4��39+o�\��X���>�a�3� c�!��Q���m�c�k�;�;��z�2!]%�e�A�dh�C���SP���䁏���܅k���'���!�M�(<�d�0Ċ1��=���o�ˑT�JE��B�Cg2|�šd-I��զ�0�5������[8}U0#>v7�&�Vm�Id_[M�e�k!&$�� �E�r�-�W�1��-T[[a��t,;�� w��j���R^*�7�7�j2Eh�j��^t~T�q!u�U�he����{�%�3s�m	\QR0���>1/b���KB�D�>�S-6d����N���gv`���9#'���m�?÷Z���z ;��J�N5bR����2�^� ��F«�@�yR)!��V����Ngw
a�(
��7rz<�dk�q�I�m��3Ɩ<������_E;�\:KX�O�ѡ�����P��FΊ��=X&�iu\nڟ�E�,<��h-mij��	=� +gJEcEAn�qJ���b�҇1$i7�<SQ�ZL&P���-jfp�Qnc���g^�H&��m�e�B%]ʲ���gqF���7\ �"����(�=�����8���^��9��}�bƞ�[D	.�q5Y�S=�~�.	Da��!�z�ZZdǶ���D�?���XlxVHYEB    91c6    13c0L�������=Y�CB\��r�"�AW��پ+�8�T��@cŽ�~�7+���E���j�x��n�����S���9+�j�>1pq�Q�f ����Cg/a���sU�U��N*�}�tT'ԝs �M�t�he1�}���lg��^z0DL����ȳ��ն��Q߼m��Fob'��#�Z�ݮ^� (&���`"P���4{��] ,ڲ2��;'kS�Ȭ8R/h o.Ԡ"��ң�����\�
S"��>�%�_�%�1�����֟d�ro�GKvl��p@�BYjDr��Y��pO��`��-L��o���v�[n.�N#���)?�:q���/�A9)����E�S`zG��d�ۮ"��OY��|?�
�4A��U�U�׆fK���g��|H&2#s�ٓS:��%=�M�e��)�k��x>Te]Q��Y>~���4���c�$$ �ŀr���-���v�����y����i��$1�P��G�5��nHJ���\H�AN��=E>`�,G�� !Ү��d*]�Oçe^0�v	���p9+Q�0hO� �2A@q�^!�/�,��m���[��&�\W�}i]\����6n���U"�c�4G�#L���I�1
wg��a(l�J�V�OAi�I�±��w�+��(��$�n>>�A�p��b�d@�Ҹ�C�׻��~�c���@�w<-;X�0=k3S�DP"R厧�K|�	��( }�s�\���Q8���y�L�y�/�� (�SvY_2FH&'f��򮷺W��H�,kߩ��b�y9V���;H�}�;:�<@�p�'�V�Q�������E)�&������������.g�٩�{��#`/s�s\OM���&k"���q��R,��@|��vO�H�^ϔQ;ݨ���yLO��~ݞY��^�X�x��c6%�Ny<@�eHa�x0W�D�H�RcDk�u��Ky���@����咺qe}a�� ��\4|���'�����Rlדk��P")1ݏ`vW�\(�@D�����`��=�I&��Z�`{���˦��`��d/鵷�i|�
BO.�!�m���~]��C���k��N�w�q=tG�hx}�
yu�1ޥ�a�
�iɝSE���z�R�������5/�wi�	�������p���̖�����ގ����tfF�zz��&]�e�>Au%��A��o��os�l�:助�Ro �Z�MU���9S��/V�8]�aD=2)N���g���d�=#]ȖO��D��֮�� �g6|n���Þ'4�5�g��fk��N�3Ro�ѰX�s}�Ṓ(#8?�Xp�1�N9�������Ȯ�����a��K�|{��J�y�CK�jz������bo�a3��?�|RWS= )�OBC���ʅ��nb�)�
ox�7	Z��1��IVǂ���3�O��7���iD�=t���;j���?2(0�vW��!����J@���_bѫ�ڦ �,7'w���J*2$`�{&�'��5�1_����
Y�x)�:W��J��ʖ`�-Ek4ST�h�Oߏ���f4���b������M�x��঵�~�Ɋ_��ET���0��6����J;��|P��wϥ�5��)!}����w�q̭*�[�\6����,��s�����U�S0l_@��w"�rK�UD��h�A�BCD��2���¤���r:��}���y�*��+�����?7(�Ŗ�i�E7͐�%��8%Q�'#(lg�U��eW}&��}��V�G'�h��OCG��̸���1�u��*Z����xo�r돗���Ԧ-��V�Y�̇��� 8��.6����^k�K[����
G
oA� (���&G��dށ�3Ӟ'��+@��9�c�'�¼��ʟ��ҽ�2�i�K�3E�s����^I�ҋA]f#k��)n�KP"� �;�׻�%*y�ʂ��/eg4V�$�����H��=O����턔0�=c�M��ӄ:D����ۑ|�	�e�\7;֝g��W��e���ti���o��=߮1a^�LE#��P���J�F+���i�~m0�V�8��+Gy�Ђ_X�%|e��|�h���sJڤ�;`�H(;mM�f�3�-���QX+R��>q2޴�`�.��N��9\�6��uּ�V^���Y���<\��ɖ���|Y��;qUȿ�2���������	�� �1wֽ�uM`t^�������yy.��`��Q㋯u�����QW:��N�3�̍2������%ݲ��{�(��j�='*Ǡ&�{�ehf*��#��lq*&,g97�\A��8�,�Eeg������D�7n���i�����|�rG�?�+|�&��d��P�׎��m�i	X��H �+��fj���^ڪ��F�3�� Ysl�@_���6VV`ƶ��aŇ)�5��D#T�Ho�����9#R���%;_�����&�|�&�0'.�D�+i��;︊�P�7�D�)2��t#4a'���Qn�`�a�����/�1�>�'�Z��N̟�^�*���UA�v�K	�coRv�&�ϭ��;�|��o�q�U�~r:��0�-�bQ�S��|���.JH����b�Q�M&,����V�R���"��B]�&aU�+���)x��l���n��o3tL��z4Q�#W�H�7�v6DЌg'Y7I�A�C%� I����ԑ������˅mޡd������yWR��o�wp�!����kjac�M�S߈�=į�&�4J¹Vd0~�r����s����4Dl��Hi0����Չ�Hq�ip�����5��bzvy��m�~o��-�!���M�����4\���ş4W�g���-M� ���sƕ�gE<�4i�AL<����5ZT��1 ��x�]\����Tg�_�^���[0�%ǋ��_���i�mtT'�)~Uj��C��"#@��8�v�!�e�ڝq%%'������]6w�=x|�ux٣u�ⵁ��Ԓ9Z9�`*Kz$�v7�J��(6�)���&��n;�W4���]+�vh\fi��hƎ���o��������KoܟH�D:r$��o}dK>!�Ƕ�U>,($	v�V~k��l/�'�p�5;����I>���V^l,��[�h!��xC����0Vvjo$�x4�葝:��@�X��wc[.Q$�ª��#�[��\^w*=�W�i3��R�@Q���fG�Y�#��#��=������$��i_m�\�_r �eg��9nʀ�l$����-Z��
x!�.x���J`1OP��1��(�C�@��R�MP&�V�f�G�
MKI �y�����%���$�M<���ŏO���Y�Fb�J} �+��"���hB�� �k@�>��z.�m{�k�K�����0&�m%� ߞ�}O��6T٢�j��wϴ
Ec�9��Yz�ՁeM9M�f��7n�|A]�����yk��W�P�^Q��=ɭd��L� �N�P��P��E�>����`�-U�q�,�(
��C/X�X���1��)��$�&�qD]d�΃�q���-jl�3�9٧� nf�cȦe�� ���OT�D2j�o.Y�+p�^Xꮅ ����H���1r���qqI�bڱ��2�(�	7���ȻN,�$j2Um9�7HN/�N�
W3�_fIG�%f�"���7�|	��k$xi�tE����.��5�������xg��$��i�5�01�iY�0���IR@w�뫸�"�)��N�+�����`$ǟGl�'��{?��B4�8O�����C�� R'���%d���r�U���:I��Y�Ԡ�1�p�o��v�w�=��H�V�B�?o��f��M��˄o��#��{�:@�0�C�������؋�W<���B��f1�=��`�D�j�z��=�"S�����b�� ����	�kT��*��;��ug�����r��n������	X1�����(.]�Qv�G�.f��fŮ��R����WYpǗK��*b�bP2���䠶8"WG�)4!�0Zϰ=���ߵ����P9<�(�z�o2��&09��З�#[�|�ͮkb��H��SO��r<O͋�DҘz.sO�쩃����A������G��y��D�-���B��I�?�n:S��d�pR��q	I�
�����]GL���GD�S�����v�t�L���ts���.�w�j�n�8�25�06�1b=�!�� �Jg�O(� _%��kE*�֯F����s啧�X��SSʦ��V+��"���uH�tNr/��g����Y�6�� F-
��ֿŹɽu#e~��i�p<y#�/�{yV�6�(x�Y\��#��j�=Ss_��IԲR��]�eSyjZTG����)�:�r�KIy�;��lմ�4�ڜF@A��m����tu�~��%8<̴�|DH�(�g����N>����
P��O�z��c���$�7��țc�6.0�0��f��~��	|g�h��j-9x �b�:�_�\Ui^kv��`T��E�dAS�p2I� ~���a��VK�yv���猐:�sa�X%<�vc�:\�04k4D@�b�}W�:��+�뵕��bFFc����%��kmĒ��I�K7��t��y���tQ�@"Ѱ�W/yf��#�O* <�x`cx����\�BA�6���̃�.��Xz����qs@ys��_4���,F
����TA����0� /c����A��bJzK`YO�>����-��h�]uoS���̕`��#��d,U�Ҋ��z���O�F�)��<�C�j��-E=�=��S_� j���s�F�����:!?VjL_�s�| ��bꯝ��{03�`	�E�)wǧ�="(���XX��U�PAX�Ӯ�r����ʶ�5:�Rb�Q�+�K~~�{}�"P*��(�ѓX>�R��,?��p���ĉ-�����i*��I�6U7ꠘ����}B��u3*�eXN�Ơ	