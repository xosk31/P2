XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����20����+�,H/���˓�%]����9}�[���6��q�k�57�Q�� jf�E�aԈ�XI �ඒ5�!B�����<ǫ60�xUa�y�J�/vCã:x��? ��/����R�^%�h�6�7�� @�(2���xH�˷�1�/^��� j�l�@��6� <~<���i�F�^��ǰč����Т�5��~�8�`gO�H&��ݡ�!�����ұnh��b��&����"`���û|G.'���vIn�Ÿd�l;@-�#{��c3��|�]�T��va&L�W��z���φ��������c����s���h�=3/���w8��ix�OP�əp� k���'�ƒ_�mv>.���}�P������2f�	�������+N{�Pk��e������X���x�PI}��T���l��G��������_�=��sD���o��V[�ZA��1r�� �ꨈ �+�������Eξ��B��_#S=���\�{bq�5��xx��*��J�
~ik������	�m�9��8�^����e}=�x韼#;j)6�-V�1�H��kg3G����@�����c�tk_w��HֽY�o/��R�2�����;��o�m��|����a����1��2�%cL��9�G�H�
��l%Ė�1�/%/��#�^Т=�8�'S�n��-�4AjJ�<㩏�/�G?���EF24x �dj��mɴ	���+um�XlxVHYEB    fa00    24c0Tul�O�6��l����_E���ltm{�n_�ؐm���~/(��-��^�*|2�?�+��rr�]ޥ��k�b'aJ,8�;�<q�7�������D�L��Dj �&çp{���	�{	nW$���N�y��0U)O �JU�؟����'�5�HW9�nB�?A'ds�V��N���@fQ�0��D8�̢��0��6��i,��WU]w�͋s��IDU�uۆ����a���2�7r �|,=�{�y�����Ԋ�����0��%-q�gם���r�,:��Ʋ�H%�J�{�漏�Msl��B]	󵰦f?��ڡ�5l�������3J�S��ߩ���_�:4��{۞��qV>A�p��dp/ %(�T/SI�j濇0X*f(X囫iFX��ߓM�%��hI�^Q��&T&L[*�ҹ��2�1/����k���@[����/8i��|�b���	̥��C�o'=�J�P3�����!�ɉh�=-�c?�hƫ�l9������/��6S���7�)�+y�G��]	Fp���3Z�b����'쉯��H�T���������B���S'�'yY�!W�^!Z��Q�j��=�^)�U��n�P�Q�THR��h�]��ōE�M�<���(���=rc�O=\�ݔ�|����^�o�	�Q`߂׳u����Q�(��î�5 O�g�~�:u���+��D�^p���[U�6fD�� �,أ��1L:pg^K�e^�d^� �T����B�˼K±�ޗ�'P!�׈_v���來қ���n�H�bU�1D#q�#IO�N�{6��ǁ&�B�}R׌O�d�|�j�)R3$�	�$��!�����j����Q�(A3с�[�ZDui��R���af?���$�&�m2�0���"dn>A��,�&q7\�X� �fI6��(8�,�xPn��^�Z�0�3�1�j7�J��p��䊾�[N�kb�jK�mӇ�b�'u\]�M�g���6����	|z
ਘL���Nå�.�eVl���SǍn��=&Vu����e�*b��aMh�a���H��� �d�r��sۢTm/�'TE�0Nj�^~֭y�kp؜4rAC����Y�6�9$�G-9�~��;0Ѷ�]��`	�z;a�m��Y\A*I�k��E޿Äk���cUg���m���Pa
��s��GD9#��m��&�j1�_��ۛȞ�`%ĳ;`�j�W�<��=^M(�5�R�8j{.��@�s7���vyo����O�Ζ;-�$��R��[�DN�7l�61�y�Wк�G�1m0SPq�Y}��P�-�.|ܑ$���%,���f,ͽSU����jR���I�������/ �ԯ�(R3���I�O��KO8�6󈘑��)$�����h��=9�j�B X7�+�����}�w��f��$���ED����1�չC<x.����F��3��B:E4^+9ٽ�:�3Z�Y\�Bq���{�FQ���R����*���ѕ&��FI�Voq��S���񕁗�CҦ�s�)�÷,���**�(cw}����)匮��B���;�^�HB|�g�sG+���8#��y��dO�$���$�5T6TQk�f�� ��4�ͬTC��U�jG2����!Ea;=���lu�����ҌW�YX����a)�G��8�����L���*�%L��2D�?�X�4� <���\����Ꟙ��P���oSDﰪ�sA=:m'9o�X��.�����A��|-?ߋ�E���CŝBԲ⊅Ȓ �;��"�l �J���9��M<�N��v�a?�a�'��A���>�  (斌ߨD��N1V���ئkND�����o�mx� ���g�=!C�/���T����B)����o�M_=җ��>��p\�H"m;h_K���sUB��b%�x�?u��dX���kEU��݃䟙� 6��:)�;%�}�����?����^�7��́lr{*�˨'���&'����3� [�0gX�I���xD2���@r��bF!P��y�`�/�=�:�����U����p��$�'��l�z��D����7�=���	�|�v��t?:�쐊��-�]�0��t|�B�z�#|aTZJ+����w���;J!���a�d��G��1�F����c��'�T�F��/���z�7����L6�d�+�"/oA';�.��j��ʎ<H�;2��������7��+K�nF��(�X�[�93Rd�:V
d�N9r˛E#AYMJ)y���=��bU����~��RX�����yFT�� d���g�9}箋S@a��S�B/;�v�gZ�lizf��=�P�8.L K��XgZ�%�'��L���y<�(8������Ť�y~��J��^�F���9\I�Ug.�����u���.{��h��EOٸ����G�p��ꗁ�_R�' �n��T9���Q�I�u��  JM�E����4Wfj�EC�ݴ4	�o��7��*��oc�H9v[Ie-g������l���Q�^�;�]�=D�M�&�._����H�`��Gi��{�6�Q14"�j�B���
��|ˎC�ɩ�&!��4@���9�>��o���M�U�r'�ԿFl�����F������T�y�o�U6أe|�|��u5�
%F'�_t:n��E�L���c'�=������Qrp؎l���O��J�;DeHl�������%���l�Gx1�� Ǜ��a����~�P�]=��*֠����Q�����
.<3tF�>�� ���L��K�m�8��� �E�~u�W���C���J`���:�(1��/ǿvί��w8��*�;*�|��Z��$l�h�StL}�6�Q�]K�'����k'V�2-.�`�#B��D��:P�H�;�q��Qj�n��\�����,��eo�[W/�Y����% ��c=���0^�թ�ٲM<��	��Z�GE��_՘*(=�Y��д�\��';}�Ri�>ո`�w{�:2"�"'A&���Xk���2���=\<��J�#ýzȓ���]���%�ΪI��`�����l����|�^Q*^��嘦\{���W��?�����!�v�֡��u���5Q�݇c8��$af߅7v+Y3��tY�?���c����~'�ܚ��%���1V��c;������
9�N%cZ���*�Q�킲P3�\ ��@��3t�A��3R�ܥ50"N�h�Q������vv�����O�rư�z�p�+n�/�t����σ�7�9W[��o<2"��PQo�}5�����Ҍ��+�7�(�k�J�P��(ѐr�G$�����Z��x��ϣM��%5�w��8�K 3wL	�
�*���Hn�k�8�{u�g�dl(�,��Y�j�N�tG˪2�F��Gmog�V�y��'na)���%�,Z~Ө����鱦˕B[g���/$����S�dN��^�~�bRd�Ђ֜8�WiZދو}�O���{���x�����x��UꗷJ[���&$�i@H�s;G�к�;$1ub��8���]?�%Z�R�K-�S�Ǐd���W�7�*���Ί5:�&���юOn�^"#
����j;q���Hc��k�Ƒ��V��C/�	��kw��$:^;Y��؞%����eת[���L�6����k�����:����1���l�'��k�ώ@�,5��z�]�aGE�|8 ���:K���5�!�^������~|ǖXDk>{�4�e��#�_�o`$�Cǃ�w���Y?�F'@WzQ�ޜ`L;|�Gt6�i�a������4�r�_Z7���YA�Ŋ�f覾wD�^�����34~Fx���s���B�$H�D�]I�t��S(��3�YpEZ~	�E�,s�<�Q�S�����G�`% ۥ���uT�U�_�<�>��D�%8��C�J��FP�Z,����ㄵ5S��nwѹ�q�^��Y��:�E��"5/�XZ�-+��e����۟�<��$��3Vw�7��g�{����[X��	&�}�=���O���ɟ���{Y:����TL�
 �&,�9��,9�	B�42|�!�\҆������{������V\ޜ<�����b��	�_��X��0i�����N�U\U�����ۻ/%���Ry���< �b	V�b�	��+럁]�	1"T��r�4��BE x����{��p��UG���-��O����^c!rd�Bx��B̥g��� +,��pq*��cĊؿ��y�J�Q2��I"6c�c����K{/�J{`���2ѢP�lL�!C����{��Ҹܕ�7F��J���:�Qn�&�Xv�%B7~��F26����6�����D���R�T�U*��V���"��Ϻ�ZK[��N�z�f�/fM��i0����ƟUj4Sa�;%�<\��D�5_�F��ad���.˕2�+X�?�������ݩdP3����WB��k3�;�F��Q��S&��x�C\E懠���$)ί�۴Т4�i�b�E^y�rcxp�_e�Z��M�/��6��"?�1|1��s��*��Tg'��Q/������/ϼ�O3e<$�G���vj���6��pg:�:�rm�p{�iE"ɳ������[2�Ů�&1FO{�L����+�K��\�����=�b�}�p���@���P2:X����j�zx!��}��
�<rAIF�+��F��)��^�8^�L�~ʣF��h��ۗC�e�Z�)FŹ^��+�ș��B`��mo�h�&k0��k,�}�K@4��W�<�Zz�<��@��_*	*,jH~�zh�2��O���r������|���r�!��X^��Lai�U��H`��us�i����eC�b`@�`S	�/�*�Ů>&�|���rr���'6[w�i���"�WY�7i���JGD�,�o��-��}�K6�I��L��jkiå���KFB�U	|���ZӜ{%�uκ�{H�
�/�A�4 ��a���=�_���<Z~C���l���܀�ߖm��޺� �����=(�=����������w��ʡk�W�4��@�-c$K���|EI֧BjQ�Z�l��J�W�U/�4���ۣ��5MG�̴��sGIL� �g�N�5I�����FƜ�\�}wd��P�*��L��qب�z�	�o�8~K��fu��F���n���4 ya�Ǒ��/3��_S��o��Q);�HmUPZ����.��G����ƈ�ݰ���ݙc��`����vn��x�.��%�w�}�H��Ί��k.�y{�G	�~F7u���LO�[�-�|_fgU��oĿ�����b[��m�
f�L�����c���F�/0c� �	�ٖ_�����WJoys�HSW�rW��W��+�~(�N*
^������_!o���?�J�an����I�t[F�S��iT	^?C��d���n����w���&�&�bp5������f%+�`w���˞z��C��(jo*�hP8��j�c�;;$tN	�o"k��F#�l��k\�PL;�'�_�LD ζ�m��f���)K�IƐ�M�_7.í���$�=���vrj�fXX^��Vĝs�h�&�E���7Ńw��u�,�c%?X�̀<���f"�fG� ��\k�L:�a��A���_��~����r������F�cB�{���Ka�ܼqQ�y6��so�D�����;t���@�@n�&��?���Y����c�%������_|8(�<i��S	�O�8�8�����QD�.��'�Ӭx�������ϯm��	���aNmZ�8P��<	&�.� {f��a!��8�9a��ѧ��B��ҩ�>�r.� C�#1����D�n@��TW}�S ,��^�r���9���l*p%=X��g�f�b6mT�e�|{����1�i7����d��\*�h���	��YU�v����_���>U7��c4|����/�YBEUX�5*:o
VB6�=;A��3�X�>^FF��E=q`���4���g%˙���ƛL�7$��!]�C���%����M'i�t@.���<�*�Ab������]kc������PP.;p����9�p����ؖ3�n�wĘ.a ����D�'j�r$���0'r0+b����r�y�1�yN���ߵȽ�ĭ���9�x� �
����P�-��l�ڙ��i�j��	�a*#���9!�p* ����aE�YF]j��+�����K�&��wo�hx�B5$bI�^��˫�9��2�\̲�l�$�_+��Z�x(0����E��Ps~)%#�.��ab=a�@��R�g�ټg�3稙�F� Y!�C -zPQ�����_O
~�pb'��C[���Zm��N�%N'�u9�h�i[��b����?� �cg�%���ܿ�a��.��΂�ʺk�8Me~�Ȋ}r�φj[�h�����TJ)���TŢ�ׅ3�a�z��{�B<.TaY"�S?YE�{����H��h��c0#����%�Q�����XQF�a����qp�C��]$�l`/_�=��ٲ�&7u�(��Y�_,)=���yq �}'�0d1�+���ջKH����1p xt��T�(�l�x:��<k	��6;I�v�3Xi� D��4�����|t�JB�3O�-���ː��R1,w�9P2�WX_�����	����:�≐θ�h�<2�ZB�KW���:���FL�H/�]ćF)�@�O}��-�eiT��(/�s>x��'�q`|�|J
�)m��?����?��
3ʃ��Rm�����5R��-2��q`��17:�Ѓ��`�<�Y�]z���qSW!\��؍Ϫ�%����%FrCԺD��׍"C� �!ԊN�d�q���"r�vƜ��"0e��A�" D�J!���f��6�V����L�Ϩ�&��I�w#�Hnč�.�p0-����F��ΜpI��߃�}��5eD���֓\�A��j .����nDW��	��ss�a�^�7?!���G��o��-|5��1z���������l���!�oOv�K-`X���9�%ֿE�L�[?��3����IJ����L7Ir>I���lw�@(���$G{�:���0�]����zJC\(0B|YJ�mҵb����e��_��HR)�7*\r�X��>�-D�&PۃBvng�ݭ��?��V�_�(���ʀ
��WEJa���ƒ�B�kXQ���m%���ͧ��4�"�@^�'X�H���\��5e�o'ڋ?.�\VS��FCUW�m��w���ΡP�+:)�R�9}���No�_`vu�3���ar�V�3�]#�$�f���IL=�%o-��Z�֏��iob9[��ظ�	�@�����:�[�O֊����jy�r���(�N���C$�5k u�-���t�E���6��b�ZC/N�,P`۝|6Z&��q�AmOuۢNG�~��{x��v���Pޝ�B-�Wްս��A�ӏA�|(�<��0����&_���st�*�Ȋx�c6���v�b��o��Jdu"濰{�c�՛�]�t;B^z���Ef�־����B��1|"��I���F�� :	�����v:o����-H�X�2$r�#�I䃙Z^����׵i����@�N�n���9�څ��)YLl�2ۛ��@�ITs}��'o�	Mͮ e�8ra��8�ɚ��؍�z y��
Qªz;��|Mw��w�g�-�:m9=�˙Ph�W)F���P����H�7��]EO����D��J�YC���Qz�;|�)���+=�["���(b���i�l�2j"b۟$�۟����a��ڑ�I<2i���ϩ�>l�����*�H<�3��7��]�b�V�?n�_�I�Q\��R����� ���4�4���=�s��q�:A1��Ii̶�I��7�y�8�r�; ������cv0�ƙ�7.J=ʽ��Y:{�ƌ�m��p�0��hA# zqi[�� Wŋ���,��A�/@�w��k��A�vT�)��`ue;�>�Q������z�s���L�L�k��J��Ԡ�N|]���A�b'VfO�p[x=�8�ŷ�E]���u�ˮ��$-K���s`a��nre���Y b�lV�S~���к�����p�1s{�,�]����.2M h��8u�wMr�z77D�u��)���4�m-.X������[����D�&��`�nh�B�郗#&��팫+8�9S�5u-��q	�N�O-	�el<�I�drɥ����z^p��.l �g��`�q����F�Y�T� �R(I��G�씴� ��F���d6��T����}�6��`�&*�$amP�� >F�˽��(�@a�9�}�^As��]Q56��JU�v�$'�Hl@���(v��b��o���G21:�2����`-�S��O�t���s�R6������~�MP�U�8���U�$ش,yF�W$�2o��L���t7s��6�	h���{PF��}#�����Q:�蜁m��C;�;��z��M˖,ZxA�osC�v�S0�'����`��h"y�`m���k]Ϥ��(��;�nۆ�݆U�����1��&��pL�0�
��:���?�6�a���f����sAC)��m����(W_0��y�����ʷ���K�_�ܻ��oF�)�ԢƄ�.�Ƨ^N�L��yڐO�kn��+i����2Uu[�����Y����S@f� <,1�?Q-Y���r�)>nq��r��i��(�X뎫���R���YNxi�E���a��/耏�<S���|D*lN�9fm�ب�H}�����QSgU����UYI�r����������++%��"R�RrBt�5z�x��vm��#t��!�{iBX�J>���_��ݟ;㥭�MJ�w�������D�j��^�-���e�����@,���@2�-�Pwu�\�t����] ��C��T�vJO���[C\��s��=��q���%��zqDǸ��[�X8�*k����,� �Di�d���� �T�G��鮠�Z1FM���v8��$�LQ����GhRj�4�¶u��ᘞ���	�$�JJ�*x��̎��	���$J���H�){�p�"tK5@�PaU�s���w9�I��$#����}�d$/V��D��|�53��C��Z�_ˠ>�dB�G��k�4�X�&�j��R��R��U�����_��/�R؀���7��ƥv�䥭�UXlxVHYEB    fa00    1e20�A���( U:cOK�E[f��	��GKY���j���Z���F��^g�R`��j�-l�N�#q�
�sSE`)����8$���6ߣ�'5����������(G?xr̭�&q�,S�^�k��bx��i��]|�y�
�h�ěhc��K0�����1��R���z�%���h�qH����fϗ>/MV���P^-���ϴmK?v(+�� Y�����dGntH�{*�(�p/z8:wXW�{D�N"��v�����t���ﵡj{���D��@�i�����.�k�5LH�8���W�)��b���q�'��	���4�'�g��}2��5��8��9�ɰPOǷG����l��TT���k���y.:t7�)�K�\��<Q6���,��qeB����J������ȥC�P���"G�G�Ӛ�Bj"�>^����#��a_mI�m��{�	��Z	��A�
��ty�˕O�n{���g�ˋZG��ϼ�ձ�q���Rt�2�<��l�����A'M�"W�]f��Sh�A1_�oVǓ1NT��ヱ�'@�1�*�(�d���v(�>z��r:�#�u�N�M��:�Dܷ���qѡ9�o�ɡ+�xu	��_P�Xx��Tǃ{[.��fx~P��Ư��Px�Ag�C�c���O ]���v�@�`uԮՙ�c`ٝ��c��9��Tz�<^v9i���R�ԄW-���8p�*�����3g�?�n��j�W��e�������u�hc-�J ʤ�����8�/,P���v���gAs� N&q����O�;�����xd��L�/���< q��o}/����F���� ���7���d��de�ݸ�]u�S�zz�^�Ԍ�?T��1/�~�*�{ B��˴�Vm[�4��G^Wx���X��U䥏�P#G2�]�t$.l�թN�S�7']`�64p(�j���?��_�,�� ��������I�<���S$�@��CW+~fzlK7�#�ѳ����<��(��"��Л����}Ahws�⭹��f����I�r��P�z ��mA��X��%���0��
�׉���cEt��@^�kV#%e���rP��`X��,>�Ò��������.��~Sg����S�]b=�vW7�.�θ}��D�y
%?d�!]���n���n�*.d�@�3:X[���9L����ĀyWH��m���������H<�]�W�p�8XJ�&(���d������S�0؎�%NW��}GY��!�7�2��P�r-������V���t;e�0>쵔e�Uw��R-X�n_D�|�@���I�F�{��R�=Ȱ
�/��l]A�Yc(x���`;]r�EɈ��#7��S�xْ�0�����~��~��l�M�ա6-i����Ƌw�>�\)n)+I�E��̒���)�4��<��(S���η+�#Q�qꖋ�Β�|5�M�v�� ����� -��x�G�/w���6������Y���C��hL*���A\�	�o ڰA�Lpt^p?:�=Yi��Ec?i���)!����j)1�%D������E����]vqZ�J؃$��;�Fde7��
��8��bg�|�b�\�se���z6q�͵�'>��^.U�\$�5',_�d�-�FXAۆ�)�I�1q̷����T㙥�M<��h���!]oV���7�������Xj�d�(���T�#IMBg�+?'E���+yzƬ(B�P�<O�a��q�VӁ���_@�
U��&�O�"�Υ��6�nM�մWe���z�b��ܨ�=��\ДI�qs��Z0��LbIM�!5ݱDČ�v̤�������	���_2ݶ���ba�O�0c���B$
<t�'B��p��M�͂)2����*"$`~e�D�TV�B�>>^xgz�i��cڗ�燮2Y�����E���q�8��2��m`ߌvagn��Kf�F(�0>��o�\ {���8$[p���d�u�����C�ˎ���
�I�@^~�>ŗ"�#ˤ��@�E6ɳ��:�=e/��Ny��/f8�W��Fw3>�xy�ZG����9�	9֥�v��-S��{}d��/d���/�t��w��ОZƨ ꢊ�כ�^�2��q�cO�i�L�^���9��Zuג5w>K��T#�� CuZ�CRf0O�§b�JE�f����9����.�����*�bgy\ǽ4�J�@p�ɴ��3������Sl���̙�i��.V���4C��7���Y۳���J����ٖs����3`�!8<٦�YM����(�۲;Ť���5���ǈ��%�ޅN�q\j��5����rD®pp=��;�a ۋť&~��i���1�Z˳`T�3�{��v��?(o˷b|�}���d��f�\���D��R8sB+��!��|&�h_7�%ځɐ�t�ja7�c��ȄZ��n�rSv }������e]eB�ׄ��͍@�zp��
�úP 5[x&Ȧp��~ 82�$�p0��r�m��y-���{m��N�k��a5i@����?��"�)%�E��)�Фh�څo炤�I�ڿ|�Byޓ!(��K�A�l��tUJ��#U�)j��_���r�w�tm�t��!�����@/ G�E�"V߃�>�KzL.�_j����q(������_[�\�����Y��6xj�aJݺ�y.R/>� $V�{�r��,|���N�z�E���I����$��ĺ���df����u�;��Ac�I/X�z��g�<��	xĒ\���|��a��g.ܼ�@���Ɲ�����Y���DW���w�e7�jb�fH�M��״R'��3J^\����ɪ����hX�ɭ�]�����l���,��A@�a���V3��)�O �n�B�<�#M�<���>�� ���[b�m����RB�I�sZ���D��@.�z�&�G������ ��62����W-!�*	�D%i�<���qh*� /r�[�5��uy� UpU�ܛ�V�˯�:�+�T��Llk{{)6X �$��x�O����c6��̷��ձ�eg�C̙�&q����_7���Ti����4� ���52�<ZGQ�>g����:�x�^�c��F����I<�b�g�"���x��V[_h�3ӯ����If_덮�qvȠ�+F�G��vZ+��gи�MK>n�w�7c���T'�K+���RN��25��g5�9��R��	�-{s����v�����4���	3�C�i��
� w�Q<�g�Ӥ��O�]��fVP����X5�1UHa��9/`��z_E��2�l�\76��@�� ��J�y�Eۧ)h"+�Ɛ4�8��,�\�^
�yS��2�ӳ!���:[qO�9�`4} 9�EI�5��{���_�[��qqX�y6�j�{�����VZ��x�B��D,0����ź{�������y��0�sO{wM`1��Ʉ^�G�������<'s4�$u�?��7��`X��W39���w�u��݃�7qE�s��n�@�J�-R�7ҎVp���������mvQ���,��������(�~�0�4q��?��*��#��ΗR�@٤�M-ȣ$�K�.����끿D����V����yH3��ϿSu���=�=��ChGR[C%�zi�PxiY�_�R3L#��V��~ʮ���>���Qrz��y�@E�Q�iH���p�1��;�\�T����i�r؍�3�^��r�B��ܽ˸0�B�\ie�s(��)��n�I���I�cMLc"�rO�Y�Z��&cz+���K�,9����ͤX����wgl� _�J�I�M��ر<S���Lj�+!囫��e�z�x�n��|1T��h����R�͖4iG��6�ʽ̻���T�Ψ���<��$4�J��ó���Q���h��_(�·��&V�;�ڎm$k֯��6���NЎwG�����~^���vQV�7�]�nL\F�G	x��2�@�� S�!UĀ9�>�� �����|���Mf?�:��1ܾG�3X^|K���Bu�7@�jNznV�C�!8 &rkV0��ZI�8O}�/�pޤ[��H;�(�<�god�P4�B��02�lTHd�a=t��O�6;�P�o%Q����*|V�^&�	]R���!���\��F
�jm��Ä/���C�\I�SO�FMTSw�9�`�s۰�l���e �4��G[I���,��6�H�b �d��X���n�F���TS�*J�%��{�D����{�Z.�!��5�y,�hۻ�b�r��gbQ����=1���T��6O�ئ� V`�?3������4\�!�|vM��s/�p�?c��N��f>�;�����
�`�x��h�����sM�2Ҧ9�.&�-?�qv��2n�*`���ITz(j�����|H$�P�������j�MլO������&�.d_����݆߹�&K�ڐF��ݭp��6���*�;O��v˚ �?�v��O%o�f�����á&t1�o��P�	���@�������0�9aJ'���g�l�<v'�D�G*��L]���D�	�O��]7~!ٖ��Wz�U���B���Re�ϤO�l�SQIE��.i&�$�}+_�b'S���cvƮF; ��k@Q�B�鸫��{7�+N>h�T�s�tZ+�8]Ta�@u��0GNۯ��8�Sa0�����s/�u���P1�p�����?�������~��*������+A/�l� �3�G��Ô�� L�sqYN�VtZw6.��Q��qRw�E���]6��A*͢����2,蹌�>"/������W���.۠ז������5(��BHYP�#�R ̻)��A�a���=����~'I[���a�L�`*|����
�{b�W���������tLѐ����%��ɥ����#@��cS����S3a�-�'��/G��-��ͳ�ng�U��Ӳ���̋��ݥQB� UL��Z��~x[�:��*�X�[|j��A���V>��>��<?�I�;(�{���Cu���0G4=���>]���$RG�S{� �6�x�$���ٽ!Oc�ɬ���I���q3��B�1�a��Zy��>�|�hu��c!KT~�t4���n�m!K�ޤ���N��/��sSwC���X�P,:�T�y.������%yDHp=JV���Z~���ﰼi0.G`�ڧ�`XF��Y>)'gt��vH��n$9�q}�omv�>��=�̜�Q���CzO0�|�sO�-4���88�!��G�n���'u�I�f���|!���E�_��ųZ&�+g0c���4��8w0���6�9�o8?��hB�D2F
I2�Kf����Wv��gnњ��颮& <WUv��ށ��@MW	�.�QQ�j��_�}i�ڑ-}���Si�=:��UR��r>��`�᭰#���������:¼s	����!�Xt^R�;�͌cAe+�&�E���T�s��0�>	?�����Qoa�!#a��!'�katu��i
c�6^����͝s�������e٤�XcA�ҡ�m����c�l�,�eɿ�$2Tl�j�~cG.<P�1�PcF-�wbY����eO�����W$M�8I�g�5�W��:��o![�^K�V�s��
�0�UmUy�u ��&z�P �z��1_0�L�X��5�V�����*�"���[�E�J�(hZE����j�`�I/~hyH������FqZbjpY�5�����(����	.���w��D�Vb-@����Dx
7DOg�C�����IhO�)��'H�a\'��i=)q�ߺ�`����G���$�RC�+�*7�so�P�C��At�,��՘�.�e�%��_�(�
����o�$J�܄�Ȋ�V(ܟ���9�Ζ)6q�Jp9���T��2Y��f|U2�:M�f/#w�9n:��^�e;�a�c!pT����ZV$;���]$��Z�|����!$�����J�����8y��9JN}.O�� R��d�����5���/OT�7�N�_?�����vK��Y�C�8Wo>������H�y�kX���[4��Ā5�JX�k�L֤����\6�y1��Ϲ2P._��/�g�b	��uvv�N\�d֏ͩJ�0�p�H�o>���U��Wg���G}14�Rh%�+�<����d�����`$����.A��8P2��8xI�v��^��������8[&��#�,� ��~�gG���2,�~#;*�:a)��136C7.������#��ތj�hn�Bȍ$v�$��+�K<~�❱6Lт�?��e��&�&{�t��P5ۋz�+-~��	���n�p��7Ɯ���|kg����.�+��	���H�;�̅���oq_�
s��Q<�l�;Ͼ2O������Q|6�%u\^P8o��^��28��B��0G�ȹ\QN��@�I.� �E,O��5?�.;I��=Q�q[����8����20�����v)��/o-"�y��^���8�:�Pd���{T��q��2m�OYO+�����,��I���<.-�{ޏ*��㺚���}�⨳���i�C�y�+J��&T�����q��F�t����S���+j,��vqF�s����͂���e��0,�vF����!�W�_���yp�Ρ[7Vm�����ٍx_�o�@�K��W� ���ҭQٺ�<&�L��.�;�0߲ܹ��_�t�ʄ���e�D,:�� �7�>R5�<��?�j=����!SI�����:!x�k6!��W:�GpCI�K�,y'�ۙ��jX�=h�U:�� �h�GY����Isagմ���b�Ɖ���٧��ͷd]�PL)x�Fgs ��­p�^�o� A�q�q8��(����^�;~�S�0�Zw��F���LX�R�EJa�����Ө�R�d�Eko`����f��~y�b��1B��A|�h��/m�a�*���_�,��!�5'
�v�����Vw\v�G���u��
`&�K����5��d@阼_$K�[=A~����'��O�@�g�ee#"vpL��-/,�,�h�0ߎ%�^"������
�3FDȸ��Ǉ�.�:,�/��ȡ��(����2���mX|W���y��w&�4�5%]-A���`u�yzJj��d�>	�,vx���	E��& _������nTӓ���`8�V����A��'Ӱ%
�t�O�2�݁Mr��1^��K=0���U�V�I��5Uq4k1#���Ur'��]=o��b{��'��d�֮5����E����1�KO������0V��'��!L���<�U*�{8y`�߱ Q�����L�3�}/N����)����e�����i8�h��P���(P�@�-P�b��H8���ܰ��$����(�~�L��9���iXt�n�X��
u)X>�2H�K�F�幑�Vy2�j�-��^���`Q( C��z�(�����8�����f��r�_}��q굚1������ʨ1�����P�"s<)��ƜXlxVHYEB    73fd    1290��
'��~8�����H�������׎��'j<��Ҧ��W�Q�ȹ�oخ�eu	j�r�����7s��Sak���\r|�-�yL��ց�AD'�m-/mL  H��&#��4��n4�RG���b�I3w)����4W��˦j!7$H)�
�ko��O������(���=�s�%[���]��r0Y�6��nrJY�����V���~�6���\��2+��)���gs�9�=�u�$���xHrGh��1]ŃT���3�UjG�J��Y3��$*@2�z׎<6*�J�`a�����k�R����\�c�F&��ր ���ަ����5����#�����%�Lk"�Q���Y	/C?��Z
��'R�$��>Z^�*��n��1<P�N
�ҽ6g@�h2V^[���>���ZH�v_wgftZ�Mxm�c�� ���}���p@#e���+�@�+"n��t�-��(�J����+�MoU�閗L!��^�� ��[�A�����H�F*��1&�5ZB4 ��C������q��ǟM3�����WkRB���Ѷ�s�갴 ��ǚ�-4�uX-���x�8�lӟ�� R*G���]h�:�ay��r|��v?i){�aۨ�G��	������|JW�=pr�i���g��e4�֭�j�ho05�F���3 ��&���d��p�`��ר�֤|�� 4M_�o�����-ā��<��sU�|�>T��v���*�����Y�II9�a(#��l��L�rg���U?Ж6J����`�m8�?1HD�q�G-y�t�(����N�v�x�k�
g?9+z���Wk�������4�
N��\�(�Ʊ�>ǕO��~�Dpf?�̈xE�1�%|���7J�LB��oSN.�!�R�]'�}�ªS���H=�q�d)S��>��["�lR�\�x�]B)�.����pp��G�=��i�t�<���kgj*u����r�=��#�]�9e$b�ޟ�*���c�sQ�d=ڽ	�����F�����w~V��j�f��֓�>��{���k[�Ao#]V"vPd/��&�-�`��zE6:�.�{fd����Gr���C}8�a-Z����q{�v~�X3���b��{��^T���t�{��nR�g����p��n,7c�C��O��p����Vb��Ɂ�T�z-��<���z��#⃿��b�o2���*�`����c�G);*�a���������ƃ��$"���D�p�5�%��)h�H�PϪ�n�����吱�\�A�i
�(�\	��'�����?�7<Hc��-%o��z�e�����3��XnEjc'j40��w9���Sm{�[W�,~��o�U���Q��
6��L� ��NIT4.x��Ѹ'��­�؎��8&��0�>�k�G?���+ℳ��:qj Θ�t��*���N�Aԫ�畒Q��fY}�4l����Dp=yGa�k�.�sz���2�j���m,�3H'|v�mZpXh�ࡖ�cUɖ4��Kk(�=���HhX%�S�.�1���k� ���V6�g�p��'�O�'�%~�(�%�D��+�#MP�9!���f$gB����Nn���[vE0Qt��d(t�0w��`���R���ꀚ:�58�������{ˑԷMx�CEN� 9��Q�糛��4�0��D�"7"�
F�L���4b�=�b�=��Rc=� <\�_��>΅`U��k�N?�;�C�`X�eUgT�ѬD�8�9�����o�<(��a�����i2V�^�����  ���+�����l��dk���!�T{���+��>ћ����C�e��.��p����50�����{-��!�)k���\�٩ZxH�QE>Y���-?�xV�I�#k+�,�sd��1K�����]Y{U~���zkXAw���9���VK,���%+�¥-�]�����x<bS���|3j�>#�4_�l/b�nzH�b�b>�����l�l�͎����NIH�'�ؽ��<��j�����oO����D���V2D�!�@d�� �W{�ë՗�[�)�*���*�I�/!���9P���u��3�l��p�SuG��SZ���ge#�^�"f�꽰-]Bl���U��@r��-�Zn�Y��\���*��r�'�e�m��S�^���[G`iփRxd�ʒr���<�+}2ȉ����/(c�s�9���%������EEdE���
3�j�*��%��f2> ��2y:������@K^�B�P���'�
~���X�= �]~��9�0���j��]ў��!����r&�NN���K��S��2�ea��B�yK:8��٤�ئ���?=���3�I^p9�%�O:���h�;����.)�+!K��o��C]5���6�w�ߖ(���!<%ܾ�����>f�+�4@w��OO t����&��܊���	/��E�����= ?)@�`�����������7�X�'$��k䙃M�����s���X����e+�|&G��mz��>k�S��O��#U2��'C��;�� �;BU�%���.�[����%�Ɠ�Ij�Z��k�)��,5���`�A�U��k�d���H�����X�o�*O��T;ɛ�˵>
������
I��x*@���;vj�"/�����λ)Xb#�� i
-Aq G��*��Kb�.6��2�6�kA�+@�@#��2�ZNl[�ŉⴕ���ܩ4*��g�y����m�$�t�BEt�O=]�!7�� YR�j�Gp��9V'��$ӄt��5s�-�M���k�(���}��y��ۻ�"(2�9�1e�Pq��C��ƻݐ�&4�ւ�gG��7�����E�Q, �YZ��o)h9ʜ���k(����� ����g�B������E�l	��c��	E�"Z15;'��'(���/,ُ��o�����*�-SNj����,+~uy�(#��R���5L�(�;!;�(�q��:���.<���i_����Qm�t�=��V�87�W�l��Pg�uA�m�FG��i��e�H%
R%o��j���jB x"q�$m){�=��R�f�=���_��t��0tgSd���T��٢��+������ԅc��{aؙ,���A�� � �|��H%�4�DM�H���꜡^�����ö*�U'��RejNC*� �q���؉�4�P���t���}�7����gS��*@7͂E�{-�Ͳ�%]���e6��=��	�̃G��N��FR�����"en�d�m,��� ^�G���u��'�.��sϾ�(�	g5�A�c������PŔ1��#����I#S�<Sĵ�r��P�x�<��4'�l
Ab|p-8��pC9���b�������fƝ�����u�b0Z�;+WF&2�+�?�՘j��n9o��xy?��t�J�v���_�t��H Bn���J�ܶ���	�t��S��o2�A�'M��6�6u��}���g�uB�ne�JJt+ W��;J��'����Bפ�aj�T� �=H��8��P���U��?�\rl�i��)��~Ttz,Ck2��ۢ��
���߹�V`W0�O�|��c&<�R��Р���[���x��!��>8�j�*�tM#÷�@��N�􍵽C|?C�%����GI�S��%B��ǴQ�,�c�f�Vm�} \��db�A~��.�05��b.L/?n��u٥=U��U,[�ժ	a�*W��jL��.�gB�J;��朽]���b¾�Po�Ή~���4D~2��|^��D�S��T�+ZH
�05�O8��+�ր�=<t_�|�ɛ��� ���w���m	e章�]`���&wSL�T_��.��r���(?>����-�����O;6�fQ�M�8q)+��Z|��ę��ޚ�ˢ�� ��"�m�(��Zw�e����{���`.=ڹG��haП����MJk5es��,nq���w���?�H�(F�s�ѩI�T����;���R-x����ɇ7え�6����>�jL��|`$������j<�!%g�`f��&�N5�J�~�0v�Kݾq�i�M�3d�A��OۯE��(g����\�����Q���wU�w��6��bS�IT�6�þ~J���\ǂ����[�5���~�o˱j��2Ȣ��=�V���[\�kE���$��l��3�F���=�֐�?h����'����yN��/��G�	���hZ��GD�J�'��D��a�����f�.dp�=AjQ�'cn3�w�-�y��sԿ��5���k;ݸ�"0{y�Œ��6uFa�n��x�ٗj��}�j�qm(�7z��+�zt-܎i���c�t���my?�K^󬼑���>�m�P��f�(��5&���#�0L�4ĥ���(�^1)�R,럭�Ï�?yUj:���7�9�r�V��"��kY�׀"	w����/°H�~���w�!Ȋ��EG{��+���Z�#���/���c��S� J�6O�?�
���[>l�<a�+ge2�uP5S��e�%��'%Ow�����x�-�������?1�(F�e����{ޚ��۝؏p�g?���YpR�pL�@Lzs��=�d`<w�u�p�()AfW[r����zy�8/���Іg����9�A��VF�JN�qN�tQ��b