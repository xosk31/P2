XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��DX�.v�I�r+��Z=��)�S�"��g��9��3&��(���S�8Xb���lR�o,�_�Z��٦�u88F���[� ���vT��=�a,ƽ�{��vZ�Ҵ����%��bE2-eV�L&���%���U,�*1�xvGB�~��A"w��f�@�����ӎ�c`��LK�g�M�6K���E��E��d;aNg�yl��OF>���0W���.�#�|��{t`w������Z�ث*�GTm�D�˘�XϠqˆ�kS�\+!��j~$�u2;ט�
@�Ϡ��"t-�����u����Z��aH}����B[��<�Y�^[�2���;�����9s�r����RI�QRL�PO�z�mn�<�3Šj�m���kBQǙ��uB,e��fS� 2>jx̼����s ��#��������od�%�&Y��P��(с軕��?_��\���*�'�y��x	�x����-���%}{�<'��H�|yޱ� ۙ�h�ݜ������ ��F
+��_��t���/ML�=_�تJ�ǎd"$�@G�����=:�����»����bH���É�����ͫ��pé�V�{F��X	y������9K�{��WS�/!#���.��0XmU -Y��[*3"ؑ��2Y�CC! _�l�QF�ċ���UʆÓ�c@�� ��e�T��ԇsҪu,at�Z�����i����͗5�p��#N���� ��� �1vHW����uH�@h��~�������N�2�Ϗ&�XlxVHYEB    fa00    1fd0�s���N?<'*,@qki`y\��J7`�.}	\�����{���E��83��k$>���6�_d��o3ޒ����<;���3F�����R�k,{��Q��O0��]�Wq��7�!��^�OZ�>	g�R+|l�f���6���oT��ީ�P�+���8$�������tG��r;�l��P����F4":BnW������X�Dp�\�XC�twJ9:���M%����lk!�' g?�����h�w���AVb�f<\!�0��'���{�`��m��tv]L1I)N�N?�'x�;90F�Yo1�ڶS�y�l@�`� �j����A����$`��������S<6�_Ȉ��w�Cl��0)X\2Lo��I'#p�P.��#[���(nߘ?KF*�k���W�j��AZ���!��Ob˞A�O6��6�P$w�5��M�&��^\���W�mM�rĕW�A��:O@�tX�b�^����\��s0�"|�����m��rUfUh��_�%�ѳ+z#E�c^ZNgpb��h
��l8σ������h����˅z�U���~剈�����ԙ�MiLY!�<��m7�N8����S`���e�;�x�Zc+�fT��hu�SF撦&�Ѯ7�Z`1�Xm�g`9�QU�U��/mk�-vZ��B
4*�����2��<v����M=�pe���E��>�#��b�q3|�0sǛ���|�^��`��)BI4�[ͥ�9g�0��c�t�1�&0	�٭��cY1��
@:����I�O����G�\ �Ŋ���-S�򙔒����	m,���-����*�Yۑ�F�z�#>.�2?�$ �<�쫯���b,E��ܟ3��qp&SbL,�AL��K����&��jP*g|.KySS�PB�CZ���zҹ�q�E"�	L��=�^:y�ǹ�i53=��ղ�Oczt��@@$��:��5�^�`�bJ��nf*�o���#��1*ý~Y�evWPݥZK/�,S��Y�2�����3іP�.��Ȯ=�[=�qE]�+V�{��cc�k����E��v\�E��ڸ����O�.>��n�X�y�s�B�d����;Wu�.\x�P�c�d���ܦ��V߂����$���ظ�kJ笽��P�6���Y������.=��\Od�+�w`������W�R���
yԼ��R�3o�
��MMb�%�ƕ�͠I��Pw ����@7�����$�,L�U��'�7��su���<�zW����'}Y�㛑)C�)EH{na ��T�\�,���
�I���<gd�h^r�ȌK�T{����<F�����G�tElU�o(L��=�c%P)z�Ǎ- V��Ӯ�r�g�9���z�vI�K���b��>�i�@���d{zg!�)?}���;���y�G3Q��.�U��z��d�Җ��뺡'��\�<C?k+�y��Al'[x_X`���_��>����R��C��S�U����N�jc.Si��64����¡���>�(L�ivˉ�����8�������ca� 4������� �%�NEr��d�u�_� b�누�����Hc�J��.��5Dt@���(��f���.���n/+a�\�*Lu'�	�M��U�I:!0�ǀP
�H�.L�ɭ�\�c�@�geM-�C`D�D�$s����It?��`�YA˥%��_ݬ3�V����9.������E���{���N?_5
���rz�̇NY!�Y�������l����s�.˾���޾����T�Y�Z�v��<� ��l��:��6wkN]g��C[�"1x������q6����.�g�5�P�lN����ljGNG�5��Н�����"\
Iv}�lV�&$��j�n�K;Z�׼-K�;&|Ǳ8-�)�Ҡ�(l���ʅ�4���Z��.J����j7��#A����$�:��!��[�:�a�+3�Vy�|��7��*Qos'�<���ہ�$��ɉo��8gm�U'����;���|��Մ��'C)_��z-��No[�ቬ	�v�U?�&��4�R�"���l��r쓍Cő����2d>��X�Q��(�"��EJ���̻�]�ҁb\�?0"���?���z����y��	��  �t���-���R� J �&�!�14�kU���QR!�}I�Y��n�+n:Z�%��?f,t;R*� ��qټh1��TSFO3���\�b�W�zN�^}����;
7-�W���#/g��S������n`� 	(��bQv��וX���������p�=.�tP�%�i�����7�]l�>,�h=+���e��8A
�t��d�j�ⷙ�	��p�8m�p>�L	��H0����TqU�b�Y`
sf<[�o9嚼�.¡"J�"�s����XJ�[��,⾩�_����������Ry��K��.��2�o���B@>X�x{��i
m#̈́�w �4��� c4�.�q�F�1B�"lN3�>�m��-;��j<���p���s�gUk1�5���B8���?9�3E�Æ朾�+�q�ԍ:u��S<t,!�m��������.��'�0���
��҄r�N���O.z%��-� �zB�C�qA\k\C�[���2�]l�5�O��	�Ι�i&��S� �Z�M{�7���M����I��ei'�n���"��3��6��E�k�&�ڑƭ0E�/�k����O�n��O�eő�&R�����7}�*�
�_�Q1ۂT:���J����Q��N�Ŀ�~�G�I'�&�	B��V���25��6�^�c6$�#�5	��.QS�솕��"�4�1_��8�Y�"����� }o;p��Ɏ��w�����d7���}_�჌�X>���m�l��#J���_�Jrߠ��֋jԾ�O ��S�`�#$�\s�)�E]�$p�m8��E�f@���z`"#�!��u��zkjx��ͰV���+����{��`���m�!ͬ��p_jh=:�}��-�Sn�3�D_,���G�z�͔��}씟����l�A�?��a��v5?#���'z�#���p�Pq��#b���B>����]�&�J� ���e"�Am���Y�&~^e��JK� �on��%�i�����tL���D�����`������栅^pH�����yE/���-N0�>N�c^ȰF�G^�#yG�?����I��V��\�.<~���'�G�n�bw[|��ѕ(�rg�+�d�r1�t�Fi�tB"O���V~2��^���j����Uh�v��3\����&�7"��n!>�3�f���t�wW�g��qj���T�R��\AzQ�"���p� s��~!2��%<������?��u��ħA��D��+�YP
�cY�9���;ʑpp���J�F!��JQ-A��Cfk��V��uѺ$�ܾt?!Q*e�ja��Ռ3��nE=$D����?�~�b8S6�Ŗ1�]k��`ۭtI����aHX���d|1�A��,�q$̅��Ů%�rK"���V��hz]�(��'��я	z-#��
np���X�����@h/�@�AB��V�m7���KtFM��P
��&�;�s�s��N�FZ}�/� B���E�.���fy���^КW��\3v<?�@��r�u�fj>��K�}�Z�%�{]���j�-B�hj������R��A���'�4�g����zu͐l�Ё��`m�6��-�WB+Mq� m���<�9��X$��E�����N��n�|��7���7r���0��c�n��i��H<�/9π㱐}�8{��Ry���q��{�^�]J��2��ł�In�v�؛K��3��}H�\���:�@g5B:�چ���Ѣ��[><�(j2Y��Qk\�	�JX��fC����p�^a�OA�b>�6�"$U��ߔ���#��ݡ�Yp�er ��!��-HUN)RUB~�rW{��M�����[�Dq��:=�]d[�4zjd ��tJ%v{�,���7��#��֫�^:�(4�ht
���NńrC�<t|�b>�)W/N)��_�Z\���|�x�$R�`��	�U�	Z�i�A�nz�+F�&��'�����Њ��v�)���2�j�Q��g���`MB�p��h,���y6�1�b��]sj��P�6'^��'x��W����?n��]�q�@�ȌM��A�+���ԑ�7:ۏG��N��9~Xd�\�/�.R�s�G3��6\B�����3'?�i���L�(0R)�6��耬#V)6�gƥ���� ����̹i� ��o����mYs�O�Y�y�-�&fZnԡ��e�I� W�z�^|gwM�F�d��Wzח���7�#\��H_�[�y+���9k\g���<+<�,�@�B3!s�Ô�w����0�Z-��9�x��xh7�����@�zJ<*�}>�;�$�_�� ݳb�<���x��^�e��hN���D�Һ�Ճ��{v`�����`,н�Ҏ�=(_��ǁ�x�9�Qa b<�RX�\���4�sQ)�5��i��������c���%��i�ԃ%��sb��ѓ!�D|�y�a�V�q�k��N� ,tj`t��nTt��ޒ e�g��c����4��'�AR�M="�E5�S�#B�,��O2Y
2�s��E�q�Џz�6��8>L�������ֈ;�=�����,>c�[Y�H�0ķ�[�z��_l�8b��pBY�_κ���31�j��������A4t�x�`�C�W,|ɂ!��WB����l����;�۠{��C"FtPG�b|����m��I��3P*�Q�穜��ﲧE��I����0��[�M�\����Mݷhݮq��kN�۠�ڵ�ᎉ4�.�4�O���`\,ZV�b�����R����������̶�T̥6���x�ʱ�����~��d�{�U8j��0��
�E�\2�DuT��,h{Jc
���m�&~G�j��XqsK�߫zm�b����cRʋB�D�ˡ]��'�ju �3���3���&v���xZה��f�'��i��/R��c��Q��#� 0�4���>�ōx�l)�4e�W�����) �'L�䱘JU�׫�w�UZ dRz<Qĥٷ����Z���W.L?f�jLs�J��p�H���&רQ2p�7��i���/��R`B�Be�����"�!O|U��cX1k�*9�4�sS�r��FW-~R���=�x��Mx���56��ڌB"��`���^g���]i&g������9V�����9p����40�1>��U�J�V�lE�J�%��!S����:B �;cG�k�b��X��32��7�SL���!lMı�:� ��F���[gٍ�������ZCGV�D�MN�gS����д��z����ЬM1�
r���r��Rh8c�3�+����k��r�%�o���JŹz˨A�_$,�P��l�c���p/O4��E�n�<�!4,o]��e9���^�U��
�;2"�̊�5xgJeݙ4�k{��3 �lE_�/l���9o2���[!�]�e� w���P�0�ַ&!@G�M��Y�H;��'�J��a�0�`��#�^H=5�u� K��*��.����k���=+^~0R��s3ӭq:�U��w��#���Op�i���A/��7��A�᩼�U=o��U�y����>�֡\S���t��C|�E��&��y���z�B����,�dر�����_��s�>�ݑ�n���ye��?\�-���!D��>�cqu�{��x��$�B�h�O������2�!�.�!l����qTHb'����6�!<>�2xDOjI[N�MG��B���G�LRk�ח��Kg�W����� ;i�0H*�%���HM��[����);!{��"�*9��z���:e�cd!��f��(y}mow %�������\Ӑ-��>�K*8͋XG��J�{fd����cv�le�d��E�� �Ty�H�
��)�T:�ֆ�od�W]Ԃ��N�V҃ivX$��y8�Ŗ��o&f�[U��m�OL��XK|+x�I'+*��S��m�-E��a�p�7$�� �F��DWTe�8PN�Ȍ�a�s��:(��)�s\��[\�N��<���h~)��n�0ͯ��vCG�{\&ǲ) ��u��=��M��&�]����hh<�@��-�Z��*3�Ռ;��cb�v~�v4&|�r�w�U��Q!��<%�n�ٸ{<�Y��KQ��Ġݸ�����e�o�n���,�I��)ş�H|���xE[@hJ7���g����o��c�q$�l�{��=1���nn����ƴ�5����ꠃp������~A�1�vŦu��|��&�֨)�^����TY�R���-����$���G�*
��<=�%`����b,:^k�]���;4�=���H����-��!�Y����gU�Y�?] qI��K�#���W�w�q�'�Xr�Ǒ_�nz;BS;��4�h�3*Ƈ�+��b�>�<�Q҉�x�V��@�n�2T���2]����4�����r׸i�}S���8���ٌD[^�+���B��X7�'2�!96;V$�{�i��C��N�X����YG�{}��nO1�D�Go�|�!q�%�˦���_��ƻ� ��RG�Ndl�ȃ�\�Jn�Ҵ�!�I���N�5�����vʟx���7�E6u�g���7�Y��L��@y���%�@�7��kə���&�B�!��k�,r Z�EeU)��/���8�:5�!�'������xY��Nդ���Hݴة4�v䖀� ��!�g�2ǩA��cc8��b� x���`��s̀�0i�>�`D�����]3_�!f2QV�Hia6a�3�X�v�&�h�^d�1 H����爞^���"�bɯ�lͶ���"��eNs_�CK?��ae$��t�=C�{F&
,�V��"/0�e?M}�=�O7���/����
��j���Z�� � G��5��H���L��N	v�%��*�
��R_u��hm�I�������r
V7����>,�
�[���(�3���{�::H�/�.=�Ǧ�I��_Pg$�hBt{�;Qw\oJ�a�m�nv���ﵽ|�h!m��mV9�Zw4:L.u?���r����"
7L�Ց���YK�Y�?#n�2���P8��B⌬EwH��c?�.��{��
��C�V������"�ahȾQ=ȽHn@�*ly�����&�@�1�=\
2��L{5��W;��`�]��-�屔��2��Z��q/�.�Ws�&��$��7*�����m	^�}����r���ҧ�E7�_���x%J��!�8(��?�Eʊ;��wY��;�8ή�3L����Iba�����]�ݪ巁�}��=���q�����x�l��	��t
� ע�[�m4˒���J"�ϝ-�x#a���̛�}=���.	2�q"{S`N��D;�g��� �!C���� ��������Nv�&�|�vU��)����M~�̻��d՟[���r�%+P���	���eu���t�����g;�#�[C��f��b��u�QIB�Ēڼ_n�ٰ�����Q��J�	�7�䡇&BS�M�� �m�p�Gf�@bU:H��\�Ǟ��ҋ&�I^�\����B�#��k���L�x ��� ���l���Vÿb}���48x��fI���
@1�⳱^���U���{u�\8��DJ��$Egi.�*)���W�`ޑ�x����t��\S��OT��3i����2׷w]����0�������@��aBKPC��F_WY3j�m�-ٔ�ڳ�ģ��
zXgV<��:���ɽ�@2�D��]F.Ǣ����
��;!~֌c��ĵ�ؕWq���6���.6Z0S���&@�&��Vg
ŒFS��N�+R�偘ڼ�51����ߺ��i�%�T|�9=�}�S�=?Bk�|���� � �x%�����s�`�.a��������Q_@,]�D�N�G�d�Tl����uO�XlxVHYEB    fa00    1340%f�O$o���^�UC��V2�u���fjg �ѓ��o��y�e�d�ژ��m�;]�J���la(r���?K��	':���RR'l����v�����V�ރмĥ�f��M�RǃV�b�f�I&�W���1,1�x��w��9����3��3��т��!� �L�L��5̫=���|����p�L���y�;�+m(�	��>�K_h�*�G-E@�Kr/�\�/�L ;f�{ztѴ�SrÄI�z9�M&�V)Ђ���t2M�?M=�����'	FK!:U��a��#��4\��o26#���h��wþ�sC�H��dm�k��I���������̌�7����2�:��GV\i�bF�kP�!ʹ#��; ��~S��0a=ꠈ��E\�������ؤ��Xz��}��D]�y�7t���N}�a:�C�{��F#��:ۥv��@�W1Kw����*IHeu<\���^�r_��� ���,͆���z�5���~'�*�̛J���f��)��-���(T�5���	�͙��T֭�!j�ޝns�'bXx3��<[5	ٟ��v��I��!9~���p���H@�!��x3 9�2��3F��9+��l�bN��Mp�~�@�i�׿��/��hv�C���:X4�Z�eYB������P䰧��r�� L���"�An�2�0nFv69�C�޵q���Z��67$9^�?U:��F��UoŮp[."�,ЕZ|�OX����tʸ��3���ɖ¬mey�F-�F�{�k��a��:yُ�&�j�c��gy=^���/��T٫�K�/�|sib�{l���2w\)�0R�Nf�	X�F�$#e¯ߟ}����B�����h[?}̒�B�N�ޥ�fJט '���0?v���%59�fB�m��v^���G��ʡ��{�j�Ylw�=��m�"@�͏W���C)����̌&.��i��G哝�qj<�
Dh�䯸��HL|�ys~���8��������p���j)Z��o�Dv�2�tb).��4I�Y/�U�1�ʰ�1�p�5���l����t�q�����Q0A!B���6h3���1#�l�J{���a���e�Q*o��P��z�E�/�GՖM�sҐ,G�X�������~3�<�,I�Ȁ�kO9v1�zcs�t_{�w�!.�E�q��������FY�`�^��p׾6��D��(>��ӹ�@%3���'1b�:y�籐~a.łW��Z��V	؟1 �c�ɥh$�wW.�y7���WR�؜�n�^��k����
�|S\S��'�{N{��&�� ��Ͼm&A�J�WS�uw;&׸╧@����Z=z�ܦhXhBvA��<r伤��_�t�)w�	��ѵA�t	�B�ɮ|��\�3�5m��?�rT��P�"BC]���e�Uѻ�'�ƹ{�����y1�B/ҥE'j�?��HD��]�(W�w��yLH���5\��1���&���E[W[V�˕�|�V�R#��s3�D��7-*�[��Z�1���]�m�.:���T�D�;Na��Y�&��'�u�Ef,��}qG�P������ǘ$<�/kiC��c������u������y�i��hZ��d�@�i	��9u�'�J�]�>��@�4��$ 2��X�zÚa�!�թG�IVnq.aa���:s��!�r�&�)uD�13o�T��|�o0�v�����1��䋫��&���W��Q��rW@�独��	u@����C�Փ��Y�a9������x�\�K8H_�۷�>Z���GF�B���o:{֯�8���}Ks���%�Xc�z���k��]�zs���{3�
&֙��C���w�����
YK��/9��Q�~*+��=�����Q��0nmq�oKdVL9>���Z�]� �5F�);V�(B-$2�&�	���g0h�8q�$�_]��6Z����[�m�3?��$�����?��N>����
���[�MLx;��c�r�E����VYr� �^�Lv�Qk�1�h�Qĺ�@ׇ�z3��x
;�G�	c�lR$[�W.QX3n�H|��pD��c|S&�Z�$�1U#h�l�tl�9��pK�޺ÝH%+z}�c�!��\�;F]��\N�w�qc�L��袊|�Oi�8{�p�r%�u!�V��cfE��v�AS.��7�Q1���FTM�凌%4~�^'
%��m��P�w���'2��6��I�D�DJ�OGۊ�s�Q���W6V�V��1I�@��0k��#�t���
~����oF�}�g�{� eE_���eZ�QrR�>�Q��w���B������UB2^[T��nX��[Z`��I<�����l��.*�-�[��3Ï����,0p�ye����:�3��e�ұ����[��JJh'*���i�g�Δ�hwe�����_��šNe���u�I�_5cm#����˨�V��[�x������<yt�����;a��W�,m��yJ�3�RM�&@�.�;�y�Z@��fw�G��;�C��E�o�����yp�s�{%��c� �<����6��P�y�������ǧ�t��d�|�nV[+2v��2�b�[O"�q �m$"��%֢5ꋮ��*��:��%a�{�L�<n;u��EE3�C��Yh32���c�:�:��{�g�x��M��}�F�"j7�O��n��^Da��ǭ���0D5ev��1- P~��]>@WT��	vA���}���f������ōߘ�/)�!�a�> r0u�\*G�U��OK��!�櫾�cP�%@���ڛM�ʎ�"���w���+cN�@ڿ�j�VݘR:=gE1��H����s�RW6��W�^w����V	=RL�\6hH�a��� ?J��<��|����o��^P+L�\��~�^F
Z�ʑ��Bp�m@� z���E�rC)�g�.��ٿ;�b�/k��G.�B�#���>pN��B���ʜ�|��r>s)5u���ZWS92mL�����)![�n��p�M�՛ ��.��huO���47�D"��1��Pj�/����T���]����Xכ+C��M���lMv�E��	#���w$(�{=��%<��ct�6�{P���<�����ɯ-}�|�V�s�����E��8a�,&X��'���N�01B�H��v-T�>��5���r�W���T|�ef{ ������e�><xz#&V`<�~Oy��1���-M1n���L>A\�N�ܬc�cw<��V��L���+D޶����a8�u����#G�=��I�1��b�?��Ngr��W ��~�Lޯ�'�U����w�Wi�B�2��h�J�`s�S��^|}��%é�٤�o�6�mxD���(�JR�v�AK��-Y�����7�jr�������G���f�9���5��ɞ�����/~��;��b^;����'qjj鳏��9�
x�^�U�S7�+�#?�G^�>���N]Z�E�k=����5���2�'T�T�ϸ�54[�$�2Y�k�ލw�G�;8&�w<�r���j?�3H��{ l%
(QL���e4SM?�� ��CЗ��}f��}�[��>&P�;�����(�*r����O$?�D(���xW��4V��4[�����z�ޔw!�HD=#�}K�R&2â����Z�< ���8�@u�V<�/��%�
�����n�2X�<��2�@kz0���S���?��;���X�k\��#��/T'�rakR��C�䐉�����k�lrZ%��q^<��s:�Y�G��ګBYC�-gT8݀RїkA0��0���oW (�b��aU�\����w\,:_>_2A�pW�� �y�����d�YI�h� �.[t��g2��Fq�ZE���B�B�J'(�Il���a��B�fH�-KF���"4�(JD_�i����ڞv������މB1�'j�����i1čִ0wtQ����0��Q��D;`ޱ�$��#<�_��t���4�������;��3]���-�[Za!�d$Nv!st
K�/)�/y6|{?w����&����+R�c�a�|<GoSW+�E�.��*m\T�!�`����*�
��ڡ��QXr��� iI�S�Qm z�ln��;�ŀ(���'���]�ǲ�f6F��8��"���:���x<��rU�&V�,��p׏1��/"רǽ�4$����jK�,� ͂W��3��*n���O	�vb!�gB�;�L9�T,JS�:4�)qf��J��uqي!�޿��
\UKf����|� ��4��������M�2S���Їf�������q�vY*#��t�8o�S"Ԧ��b��]�ȷ7��6Yz�Y}��#���i�<}�!���
��AS}4��A�n��z�N�mj���ҳ3��-Ѭ������9��ͩ���ef��U�R���`���Wl2�L�=-4���5Jߡ��3��g���\��K��D'E��.��8��ٳh��^:�i��+�PcPۄ�Yʕ�0L&�<&��~Xj>�8��	e${[��]4�`K
�����}I�������j���ĝz3if�����\��`�m�t��w۷i��c"�|6���[*�4�<�O���u���hM����I��U_�<���D)��|�왕�#�_P�����>�I��TK��5��Z�Gi��jl����- fcDDX�	oO����ɿ1��,�O�WO���m�-I����h�&����t�"q)�޸���m��Q�K<̦+k��ɘiw���󋇫��[��J�l��
N̲P�Żx曯C�#��1���Z��N�O��{h�Y�Iƙ�h��9�gH�Z���"�83�5��`|	tۥDC���XlxVHYEB      e7      a0v�5�<}���-���T|&#vP�$m��M]�6q��ܽ̃LУLi��Nov+*Al�i����*c�8P�q1�z6F�l\�٩���.SZGz�=�:�^��%Yq�91y4���p��� -UXz$@���D3'�mg&
�	è)��+t�_]b��[->k�#ן