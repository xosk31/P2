XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���$�5�d��XE�tm��mh'��KL*}`Yk��k���+�j��y����Dzd_fk�D��'	�L�<�|�-M�5N��5p�*[�P�Ī�tzD��%�A��,�'�0��`�M���[ ���ۅ%=g�l���	�}
ֻ%K:���������d�"ɫt����[�ɻx�h�R��6Ɨ���q}���R�)2�s���W;~/���/^빟x�����IҰB��]��>)Pأ&�yls��1���R_ْ�d�O��ۮS���Kz�K��5�H�f���V���-y�>:;5��T��P�O���2�K�8�4E��A׆(�.=M׭�ozﳜ�s��ܑ��6���4�����Xݸ���*�~�2��TO��Lƭ��k����R�7����C
-��A-Md���Ŵ��$��{�.�Cvo�����i�m�Q��hX�,@�C:�&��h|i���c�$� ���6Ֆ�����c	���z��ѵ��F�iQ�����R��u�#`��6=e�I���M�f�J���f��MUsx&�{�&p��?N�ͼ�����]�m���18�����5�#��8 �c�O ��~�c��`|��EVK��S�����7�Oe�n���3.�#ۋQ�����`�����	MV�u\�q��F1��i�
W�_g�7�ѼG�x��a6b�De��Ĺ&Ys�z��~)lyT����U��4��� ��Pj2���:�T���Dr��۾s�9�%���n_�;�n�-XlxVHYEB    838b    1770j����0��Ì?�h�W���?\`��|�:G=�Zr	��qm^��m���c�X��,�>E˺ʠWXJk��81Wp�"���=$Mm��{�PO (s�3_L����"�`f�	�z7�:�[��zMT��`I�.Ms�"��l�6�:;���7��p(g�����}��ҡ�^dH��ׄ���e��C�8e��Ĉ��-���Sӵ}P"��@�[Q��L3��RP����%���((�#��c�'��NN���CibɤSܖd��Ow�*W-n�v�P�j��=�'p��f���Ru���e��г�z1ȢvxE�8,Λ���Ф���T������h��(N���pY914�\ �{��+��5�����/I��^s�σ\���G:������j �|�Q)���V��N֖r��0�Y���o5����l-Tk�+��&D�s��3�W��
7iX���R��k�J�G1ɞB�[��N��U��}��Tg��(��@ަ���$
��^��� 3���Δh9�Jo�9g�6�oc�C)�r�e�X-����Eo������EV������DE�&��
1��]�?ɵ��pnڸ�(	fY�����	v�28����N�F�r�#\9@�t��Ot";��P�G�����1��aY�jh����|�=������ -'�pR��!����L���m�Y�`cSϭbq�s��q)���x�В�*n�[a���l���������
f�G<�>]fJ���x�z��NOr����-�R!�4Y�1'ϡ�{��ZCɆ����G�j��)�3�H֮�;�/b������#)^3��=o����A/"�|�5��H�X?��[�|���'ބ�]�l�sM=�u��(%?n�%1�����y$�ue%m�91)�Y�l�
�O[v`K�z��U�,O$�BC���a:���S��{{۳��(�C=���
��EX�Me����tRF����j'x%���sH�)�?- ��$���S��@��!�,8����	��tÚwR�c/X#�iVɵtH�oǙ3�g��#(v��r��-B��&K�iO1�w�N��j�-?�����x��(�+%S��&a/q��2�+�Y��;k;�>;�??��؝&�}���	h}Ć��e���OqGcڱA�:��33�����A�u>@u��1���O���I]��rՔ��ƬJ���,W�^$�5�y�Cѭ�v��-)P�C�G����/0�]�J�@Ixsa�-`�z*��F��Οf1�H��h�X����L�@�������Ϧa����ml���Ύu,:��Y��c)q����゗�ڟR�y�-��4f��ێNS���3��0���`[U-��������S[K&����J��32� �$]���6��)�U��Y����&^0;?b�	���	h�m��w�Q�R7��fq�����|\d;�&�@8�BB�x�(��}z𺌊��n�o�bp��᳷f��꾽���_U?}6��2�L�����Ĭ���� ˥��t����#f��a��>��C��M�>v�~��+������[v���.��WЙ��W�C�n�w?���^6H����y�(1�&G�+��+�H���á�c���tJPK����2|Y�{�K�
��g2�Dn�	]����S��&g��M��t��2��ߠ6,��E�C�Ji�[ƕo"�h: �
sB��&YNEOgH� ��e���0�-��.�c�M�Ь�YS���?�W��̚\�)Ik�B@��=��� ��nڐ�-ؒ��u	���u�KAiT����@ͯB�"��22���v���	fT�q~�p�f�R���6+L ^p"TZ�H�BW�+J`�MJ��U��\2Ϳy9N�H�M%��gf�jʥ���k���X�7��j�3�s��W�u{��XP3�ޞ�����|�q�xe��ǃF�xjaY2_;;	r�"6�U�x�|��C�ۭ~3������,��&��ٷ?�;Kü���,2��ert�����c�9]
�.�G������,��Y➧���n��A	��<*,�-6��������|S1�{����bҌ��Ou,)���H\ӮV}�_(�.ߘYK~?޾p{��,�*�C�"����"�i�c����t��h	y �{%�߾�����g�G���W�8L	o�� �a��e�������� sE�~x��R�ة3�ȿ�s��pH�HZ`�@���	D3v'�RuZC�_�;��&�y�M�Պ�I��{8�����l@A�"R�R����!���nK��Mj>�w )Zq�igH�ӄ�oai76Al���'�u���Ŝxa�̼�Q�Iqig�uj�g�\��*�1�%,ћ��%Y�q��Fa��_to�d�/��
�MA��������y��&A�+�G&�^��S�N�ͷ4i�GsUE/��tm��*�t�J�ԛ��7�1��D!|���-J��?�J&g@p���<t{������h�E���[�(�Zk������vk������d^�h9�y0�E�B�L�\�6�t�N?1�^{�'G�=p냺�A�?5Q�\1=޵�Q���0'�2�M��F���TOq�/n��*C�D�s��[H�a0�Fe�s��2�з˕'�S��{ޖE?��sQn�"����R§/D/�_��!��^�x�!�,��_�h{����;�c�6�Q(=\;b��b VB���o��>o]>�[��mq��}��C��kE)՚g_{?��A���;IM�R�K���@W�qC}m}f9���]��*!ˢ�F�IC9��Hk/x���z��;�i��(���G���*J��R7i�KE?8�e��w�M�����x��ـ�";���X�^�S"E��q$
+��z�%|�J[j'(&��pD%�JTn�:[Ds����MX���5�)np�Ц�\�����b��,����6�����|��	�2�����
��\񏅛Fj�꟥ml
��:9�]4�ccG����~!t�Q Aw<�m�� }"~+����1L���-�`�R��ɼ7#~P�a(�wf[�Ս|��4� ����8o&H���u����X�<3l�C���~�OG�v�q�ń��6���a��}�%��mCz������E��"C^W��\OMW�~�.����N1FĤA��hX�uS���gg�����B7	�V���k� Խ��}B_� M�SE�L�Y���eX�dB䋂VȎ㸻Ա"$�I>�Sme��s�j�F2_��-��a��;Ūw�j����D�◽�sR��Rču��\���}FPז��X �:��>��x5MjrG#<�lI���~�[4ө*dV���twL�"o�G^E�ϼ��ƾgt�猯9�Ɉ�V8�x�z�޻�ݓ]f��N��a.R��1�@�p�Ѭ�A[��Gp�)�ϙrk�@=L^g�{��xs�F+� ��kh�3"��M�uՎ$��@���im�ػcMY�%�]t�b�&�ـ�����������7v�Z5lf��e���q�"�/��m��2C_UD�Z%P�����y�V��K�@�R����VaEɐT�{P�`�mz'�7o5t���t�D=���c9ZB�L�s��F7�~Jq�ŋ��� �L����l���*�F�v��1�٤���.H;P|C7�/�z�8��A����3���8��w����L#���o���X+_k� �4��C��HȂ��E�-޾<�MC����`��J�ҿ&������UIY ����Z�?*��9���v'�,�u_�� g�!�,@����C-��$e,��dq 0���8��륦�V������=`TP8B��u�j���H�\���͔�C��*x� iT�,x�& ��	�lR?���B��#U+f���&�7�&fn ��ȸf���j�B�-�=���ؾ�ي��͟q�(
�(�����0E,ya���q�]�~�]����K�끫q��"�@G� M��YP
�����i�kk���1�,��qtߺ���n�|�,g�_���EޓF(t�ɴ|�/Kw����Ȇ�1��棎w�����ԝ�|^0��IP���0�����Z`:A�&�'�cdc�N�;�u��zQ&�k/ʍ�G��㵈
p[�,�V�*ڍ�t:�Z^٢�Rd��ɞ�V���/��e7����< ��ڣ��Fe�|NN/�]X��1J�S��nƶO���ET"w�;��\UA}ނۺ-��A�[I[����'���ę4C�pȧ;�W��r/o�G_;
�z	�Vz�RA/7��4ҕ����9�7���7Q�񣓟.6m7-�����O�׳�`��K� �<��&�N����+�a�Fk� �s�a��#2��l%�FVe#[��-2�h\|�[n��0]��vo�W�ӎ������Я�^���Im���*�����'��8cq�"��[�P����"�6����2�Ե��%� �GUl31,�Za����Vݡ�~�6��CS�d�G��)Ϋ�a�\o�X=9/B����V <Wy>./v@�P�t.$��#�[����QPu�/��	@��DT���OqכTDr�š�L@���������'�2�k��]�>~l�<
	��x��� �/^��tG�@Z�#�<1G��>L�p�e����$���,�P%����_7 e�/Æ�׏��k{H>�h/y�{�I��@�i�M���؀���0�]����88X���KŅ�5<b�Q}�^�7�	V7:�0�\����uoo�;R���"�P����O�;֞:���m䱎V��,� �K�7��x1�� �*nʪ�ũxEgֳ'�*��m�\1 4�%�>f�Ka�Cna��xп��C�R��P������R-�B�w"�0�~�Q�����=��+�
}R��p��^�9i���Mb�h�^���M��9�GS��+��'S�Cㄤ�^���a�s���I�%wLG���nA�V5�>N���kQV$���/�6,�/c�����Tu
���)�#<)Ί�uS^pv�Nj�l"��U�+��_�k�W�c��fc�ֺ�]�u!Kˁ)E�^��:?��
?��Nx��&������dT�U!zk��,���Cn�|X��p������$V]`!�Nd֛t�����Tւ�N ?K�����n�`У��J�P�#�Ml)�t�qe�������K��ґ='W�x���!&p�cX9V�K��qZ�>#^ݹ�=�����K}�K$42��䩌���05��G;�K���Ad�"����E��"X���#��d0K���A[�<}��8�)V��~�bQ���6*�����ԩ�:tX8úҤ�qIrX�t������PwݦD�0��N$�ҮȂ�*U(�[ܲ��^�6�/4��g�Dbf}mD�����$����v$�a�K��ظo|��Ly������շ!sY/��E:ð5�t�}zd�b&����vu$��ݴ,h?�j^]�����Ieʦ�EV��*�����~o�D�h��YƸ�
r���$[�;4,js�T.<�7���@ƀ��+�^��{3j�_����i��ݡ�(@��ݣ���Yw���[Sd�sYT��7X�Z����O��_����Ֆ8{Yb�޷��c�}3Gm�uS�\ \!�H�/K R!F��V�8�T ���'��e��D/�������jle�9V�`)O�qc�u)� ��+������i��5�&f�ͧ�y��Y��֟r�g�����z��������W���p��k֦(���ʔ/��mM�)n6�-��7L����v�2�q`�Xc�(������ߙ�a�I@��	הf���ѮU�,����8�LmD�I��h3��Cs��ua~�5