XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���c)��w��7�k?ɷmLJ�|���ߪ�Q�9���� ���/ �C����ZxB�yJ?�,�66�3�z~�T�S�A?U�Ea<D
����L��zH��F{�D�T»��SG��2;��>�;�����,���(� ����jYu���H�"��~7�ؾ[N�� Hm�nl��!��a^y�!%�6�W?�Z�a:s�\_H�`֨�����-��6)@O���@�_�!��]ϧS�(�fP~żB�6=H�,O���O�o�H<:�N,�1��;q{�`�)�w=�u����SE���Y��	eʁ=.�	[�#��o`�%�Q9%]����.^��=���
(ܺ�C]V�ݬh֪+~uɤ)-�F'Wc'	�ɀ^B��ԛ����'�VM/Nq��b��f�N���a��/�_��ș�b��^O�u�Ҧ�Z�ޚ^�b)K�֖����r#��Y�"��W�p����n%w�0�G$�,l��ӏ��ߦt�	"T_W�|�HM	�&^i{'���V�x8p8yO�9P�V�ե��d�vn�8^W.��4J��� #�V���1B+/�����bt��F�B����4f򣪉#�X^�a�a��<�#˿�kiokK��%t~R\��8�*n�0�쫳��gQ��GZ�'��M��(��vr�$o���U�6�Q$�ˆ��4�Zph������}x�yN�Ŋu<��d�=B7L��b�A�QP��L/6��Z��gK�3�x���]���WV��o�QXlxVHYEB    1ffe     9b0������w-������O��r{p�v���˵���`EK yB"���^�9�@���ԺL+�^��=zҡBs�ɋm;��h�$i�� ��a�s^d��7�VR{��Ʊ�	�:ɛ͜�E�i/��\�bm�\bɘ��s����ɮ����M�b|�؏�+[#�~�K�m��7g��P%�%o�p�38�}>$<O@"0@�U7-UF���J>��rM����[i�H葮���ŭ
��l<��w(ă�j�&��ʡh�L���G���&��'{G^4���O&��a���h'r��2�iF.st3W�S��_Nŝ.���^�K@�Y�\�s�/��9f������ŰYDÆ������{ӓL�c����G:/�s��pS��dJ����|pX�c�@	/�4�b�Cf:9�@門x���xO�;0�\�!yb�xq=fb�
��|�&�T8�5h�K�-X���"�d�Z� %)�Q��(�Jf�������NB������ͳ����i�%s �MN����o�W�����x���U6�,��y�-)�y��)RKQ�nRh�_HQ�g>Z���~Cà�ɸ؝�
��o���#S�b�`�T6��E-utwԺ�3MO�1��3�WH��7s�x�����>�8�n
���������拉G��=E-Ǹ(��dii���q`dvf���O�.�}�Y�q�o�Vw)�9{dʍ�Q�����2%z;��M;����T��,e����L��#Sb_�.��(uz�6��>�~���2
�Ǥ5�eJ8�����zp��K���F��<���'�?0�k���bU���_���<t^���j�H��g#�r6�X�.���bM��ѣ���˨{���X��l�i�X~����h�A�ۘj�QO@�enRo^�����j��Y�*0%�8�}uʛۨHH�R`�q���p�r疄V3)Ki尷%�ؒR5����\;���PI��k~��#��@
=��M�vԆUJ��H"'�>��|��4ľ5�iz�o�; �ZTmjA)dx��1]���7�����z��������z��DVO��a���4��p��+&2e���J�)m�
R��U���o���Z��Şj��=m�$�]!#�!���t����P�@����`�<Gd�T��9hX�4�jp��v/0�C��y������7��nҏA;O�L��M�ϰ����R;�U����U��������w�eK�^��)a	y����Y��Nq�O�^r�N��T�]�E$�\�|'�`S���A�c���Ȟ����`��]f^qW*h�"�TV�-�����A���^#��A�'3Ɩk2+x<j�G	��vVaER��y���.�x&׾�nuD��ť���]R����)����Ǳ�S-^���b����O��{Z� B��5'T!(JQ6�k8GkA�C! �%2k��8����J��Ǒ<<��Z�/gqFN�q��Wi'�;S���BY�>�а�$�P>��^���^��O>�j���r�4������U��%S�f�;X�d��p�e�)��BL�H�q҆��c1?�˨c�Q>ʫ�.d�9��7��K�HEdk���4S\�,�G��;e#KA�{��O~&g�k@l�6����`�-�i>� �4i��U.A�?�5ޚ�)�~3�g�Z�w�>g��?�<����r��.�ܚɊ��Կ������v�8�1`L��5|b��=��g%![�v�c&�#h�S=$��y1tr�4��{$�݀4 ��lz�>k��yEP� V�{ֵ@ad����;������B��U��@w�d�
��)�# ���$����h#Z��������y��?��_�Jw��x�6r�"��_=?N�?���� �k# _z�D�5f#����|��!f���� �����{a��L<�x��J���83q���N�'�N;�w��/ʉQ@�nm�P?��w���6��L��.�¬�W�焀�<��/��,|o{��a^I"��ܑ�
�H ���&��`z�����Qӧ��q�!u����BE"-�/%=E�Ă��_�����֝��Fc�HW��o�?�
%�C��/P�{8���0�k��c(1������,5T��ќW�f/K�{�
�������V�k�<S{����*��-��"��|v�)[y(N9P�\܋� �7<(3p[�����l0��!��^��.�\vJ�$���#��L/�B\�4�̆ݾ���F��5���h>]D2��Z�q�� %�������G�<��^4ixWH�T�<�Z���ȿip� �L�[CΆ�����nK��I��$��{Z�R�b{���T\^9ރ[���^8�����]��J��C�BN��=VME��mT��v����lϛa��g=�����y;c�9�!�#��?G3���:�(�\����|:C��R����<� ��nW�7} �N�