XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ߔ�k�&��B3��fu.�B���l����S3��X��E殕"+=M\��3�����IۅDB�p���Z�C���kJ]ľW�d��Q�Q8��Cf��0}��{@9�y8 k���9'���R�Z���\�J�,�/T��@ʢ(�V����_�:��O�+���w����p`�7�#���(��h���Ԋ@Ο$]"����"��V�K���*br��f��{h-k��T0��L�	�ބW��C�QI��,}�޷i~�
]�E�wf�� ����Qk�Ǜ���H��ͦd�����ғQ�쓕r�.���[���Vze���j���|IȀ�R;Y�Zp����O��r��hEuf�t{�m����3/Y���D�7( �$��n���sVg��#�Q�XK�h� 蠷��#��$�J�"��[]O��/�!��Mg� �;��3�b1����J�Z��'���|�u4�mG�q>D rt}!,>��xQ�r��/��d�	�9*~xs {�6����w5,a5����]��z�6�V�iBoZ,�7g8_ȵD/���.�p ��W�I�hmZrv�C��=�b��Ƥ��l`��j1�z��\���؀ʪ�^��ѳǉ|{�v�8ս]E@��U��(L��s��XC�L<Q��3�d�^&��}��v}��4 !�e���tw�m�HD�o� E�H�y�塀19�$��C�Dt�b�7�W���t�<�D|@����v?�/;�N� ��ʾFXlxVHYEB    50f8    1010���C�%�!a�iȢM��Jp�#ǩ���B�h��3�U`!^�ӗ5���=�3�_��S��"������nC��'s�)�ݨ(�$겪����c�@����Uh����[���<��G��1�)nr��) �t��D5"�h	H�q�T�9�?.Rt���l�:aeIv!4�*����E9�b��{If{9 �����E���je;L7r:�O&Վ����_��c���)�i)���>�>l���� i��.+nP?�;Dk�������r�U�/��v�4iɰ*�T�%��S��5<ir�v薥�Qb�C_�'v._��Jr��O�S����y~f�;��	?���!P�;/v���W=7ѩn�c���vwcRg�@����|j�[ϒj�7R�]�^)�DL���zn+�p��T�b bi�&�<�Ε�TM���M�^S����ԫN��A�_
��˕��'� �Cשּas:aqn��"m(Z���}�v�,�X��D*���B�L���i��53�^�A��ĥ��(�1��q���(�k��^4��5�������%����T�#`�R�qś��X9]��NƗ��/�GܠͫF�R�e.D���`�I���D������7d-k��Q�.��Ȝ�i7���$�9F�f��6Nx�y]�!��
�sS?�I�Sa�v3H�!��cfI��3���"�s.�i#;e�)ݸ�M��'dބ��y��+�����`�,����E�PH��/�3\�mfV�&��+���R'���֕����!�O�Z�9�fQ2w�r��
�B�&\�j�= l��Yp%h����n����#��+Zgao��0���T���W���h첞d�u(�휡{tt
�^I��w�ztV�S����=#2�"$�_���=x"��V�u�~���۴����Wp�&����0Qvo���훴�M��7t��@�	L�5+��(����~�rW�O�zZ#_w�����U�m�����s��oQ�?Y_�3���&{���N�-�P��n̨Sr�Za+��b'!��u�<���rN�S��ِ��t��<�q�P�/�Q�-���)����'������2T�wϸ��V�gx��Qٿ�B�2�]�Fx	mn6i��8S&���}j�_F�2݋�Ď�]�C�������T.���1��K��TZ�s��[�I(�p|غ@stl}ktbrmg����g�#��#u��2�����; ���$�]����[���Z-�D�*��&O��=��+�qƗQOq%�k�����
8ʃ7��}܁�b?up�_v���-� ��ه0�|۞Q�c<
U}�'W�LE1�ep�|�����n��|+]���SY՗��c5��
�S�Xpx�$VY}�D�gޞH�h���������~�6�7T^��$�������k�5�*���ɾ�v�� @�����p��H��=�qo�( t���6�5ɑ�D �f��}KeT俕Қ�˱��gz��1go�2���0���i�ko�?z����ti��Ή>����'��l���d͞�5�L�j�źY0 �th2J��{I�%U�=[��M�5d ��͡��1���C1��2`<F�! {~v �y"����>�����j{l�b_�֏#g���t0�:i���I�V"�ز���CT��P7S�گ�A�D&$���b�Pu-ҕ̛}qs�_:�\�J~@4E2ý����A��F˓�LL(8H�kq�������{�������a�R���NxU?�^���2j�)J���sp�қ������*�5���hx�ۼhG��*��G���3�XJ�{���W��3wB��J�W�¥=i��t���D��!�N|��d��O��`/za6��kL�����j`�BK-��,W�Ny���v'� �H��\�u��X�{��Ӄ��nV���I������i�tPR��B��m���.n����TJU�R���W�18�9�D_%Ǚ��ʰ><�bY(Uk��h>��Rܞz�PY
��X�((�=î�ё����?g�ol�%�j�?�	d漈q;��l�Ɲ�#��&���T�O'��2i���H�4�ތ��ٸ��u�"���?����S�X8-�?ތ#�?�J�x�=��O����
U7>��d�S��H^2\�8�^VYG"o�%�:hp�E'�����V��\C�1���C�H�Z/�s,8��-u'��Uy@���Q;�;]�p<����������-5�̔4T�n��v?��TSx��^�YV��[������bGT$Er����s�����4v���bNΨs~�3�/c^����B�=�[��5Ӥ	��Y���{��ۊ�����%F/�M�2���ܾ� ��b-EDOqc�����@׉��	�iJ��H�'&D�9�x�%��>�Z�%v���K����Ѿ��ύyPd��vN5K:��w���G� ��D1����4�|�E@�ԭ&������$�J�.}�R����J$܁����W0g!W�����z��d������/Ss�&��u�J�KLb�0��NG~R{�r�-Ö��}P���OaN~���f�����;�e��!0P5�/���)����%⸶�ڧt�t��EB�wݹܸ��0@]
�I�ǁ&".�:���2�/�VJ5{h��fm-�W��*͑q��5֥�0��{���~�>ٵJ��K�giZ�$�*ܥr�aG�J��8����V9˫�>�X�W�]&�ir! Ӿ�h�C�(�i�y;��}頮�Y[O*t���	��S���Nn T�;�2ŞG���^�:�2�:������;���h(j�B/�v�+�����^]0�zD~6����9O<0����g`[�I�k,�O�H�Y��r�C��#V�U���
|�W����Cf�q�r���X� ��Ȼףv�]���d'����������~�ؿ̯��l�M����A�rA!^	���
����]�-/>f]�
rcjF�In�M֫b�l���>��X�+�W�di M�H��gqj �h���vΡ[e����M�h"m�E�%fؐl�4��{l~�F{��5�D>�l�1��י�lz��p��ir�RN��O1ȑ�2Ě���t��+�����S9�uEc��C��,#U\#�B�I|i�L1��FiN٣�0XM�����s����qӖA��}�$�ɞU����/1����0��P��O��NK_N��I_lwrDm}���������H��.�7,�R�]��ֆ���	
�v*B�<��܅�Vݼ�y=��9]qR��sR)<�����챆�~&	�$ӚG������Cl��6���@T�'rXN4��:��>�L���I�S��Am��ak���P�SGq1eQ�^�M�P�3���V?����=ڮb�4����,aD!������;�ډ,ձ��'4>���^V��H�>�G�q��4#K��o�K��4��82I"'ڧd�h�+So�Y�(�:���]�ei�)��m���:��� �?�a_pY���&�<R9-�	���,��	�������E�ࡓ��c2�a��K,p�0�¢����#�{Q���T|hZ#uZ=�b%Gt�r`\,�~Y��A�cpSrf�S1vGV7�A8j���SJ�`�h8J;��z�D�7�"\���ԧ݌�fj�Ί��Zk��ڸ���+�X�
^�&B�Fٞ�9�KC�����Vmm�� /�=o�/�9���� �9@Ҏ�K��)D��*�	&��j6 ��^���}V�Gj骒tC@!��l�=9�2��z;iU���
s9���
�}ڐ��rtқU��Z��������R[��d�A0��Y+���پ�	�՛�PE�J����;�6p�?��3=����'wx�;���}�F�'Rf;s�>�q����)<�v����3ps�����'%n�)WB �E�R~l�e�`n��ɷ`HڑU!Wrrb�ܹ�K���;�l5��{��,��������L�L1�u�i8e)��	|0t�Id�%뎔��x�)6������s