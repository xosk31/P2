XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���aiwISP9��7��ѻ��q���z��ᓅ��Z���(�wo�=�C�ʧ	�ZfK�2�l�i�	��y���jY�9�	v�a\����s���5�>⊵9
��+S������֔�^��w�X�ݓV��A�WY}��;RHM��IOas;��K��ڑ'ݿ�v�F��ě���(��	pY{�P�%Wf�2�ϸ���ԍ��)��%�*�ʯ�p�8+���'j�hp�?!M�wO[X$C�wUM�P�q�!	ڪatbG�� p7�)y�<��[����	�o�6��v��1ۈ*�؝��"�YRV�;X�`��r��󝡽դ�{L����\a�`<���M���!�j 
Q�|��bN0�����?4.�ܴ� ��G^Ԁ�I��c^����G<�H!u��Ig��m����k��>�|x�_��Ǽ6$/?ðR�y�06��f�L>�
v~��\����ϰ�ح�j-$Wm���/p�x�V����t�r~�������Ȗ������8��Y�T�������7��4�r��*�}T�i��Yg7�'�f��W"[��N��	{�ilr̡���i��9H�/l���Y�f,�'(�>uhp
��-����%'�1I�"�,����m�m�Fz����-RR���/(|O7�ԣ�.�W?DP��5v����U���g�q)G�3�D)��a��>��v�rR����|��XK��Z�ʰj���f@�R:0hHr�J��*�R[#�4�7��Q�o�XO,�l��XlxVHYEB    130e     7a0j��^��*9b��.��[A�Wj-�Q�S�Ϗ�wY�z�+���Y�-+�M{|�;�s��#�H���O�m<���^���zsj�LT#��!�s�m$�H��ޠG��]}槃�����i#�\hU�U!3��w�ڶd>��x�n:�j��dFӐ˱�[oR�G�S@$i^"���(�>;�s�O��1� u����c�˘�� ������D�[�+X�PqOe:OJP9�e�Z:ڣl�b�Lg�k��n��^G�Z��s�?n��B,��������h�7�Ʈ�B.F�o�X�5�8L_���=�f��a���F�t�����Bl�=�H
"�:� �M'N�9��}�1m崔�~��ʞ�P�j���}e���g������(U�bsd��N(�k��C�r�z��R��7��"��|�d$�|X��6��j�0x�����G��w0`�㢊�d�XDM���i��:�3/LE�O�;iH�N��C7I��H�H�S�yO\��ܐx�,.:�f��Gg�1ܣ�̹C���L*�0m��H/kP�.��Qi`�{�U��f�}��9d(kmH�dO��G�4;o�?�M�r��e!9]��E���]}u�mwJ�6��%�l:`B��Bv��������2���!SV��8�w��C��@� 3ny���
��,#�4d�]u�+��r�����\=�^��y\��� ���/����@�.�C�:�jNv�cmc��n��)[szSM4_sn������y�[ދ�Kb��Z?�
�K�7��MޏY&��:Vok���yRs>��K= �JE8
m�B��jkfb������ ���@H9dZjc2}�
�]�͠s�]�
�x/��
����M��KJ]�����h3�RKX�x9����e(�c�9 �̵����r����i����փ,v��N�rSl-������nL[���L�v�"w�����z�,;���ڷ�P����֯�I ����Q-�9���v	y\�U��ߟ�oOU`��~|�9����7���y��I���,X�����1��J���!�6��ْ��yq�n�4���9��#e5i� ×	����v�"�_ӈ��8=%,=j�~���M�1iI�]�T��8<\%��pkƅ���d���ܰ���D�X�w��$j��.5�'�27��W�2�q��Ȋ�����5"�x1�*c�^�j(-�$%��j
aI�!��H�"%�o@9=	d����鯈�'50������DTj�}�J,��ɕ:�Y�?Q4ҍ��������T��o��v��*���\_TNG�3�����ga�!���\�!H���t����$���t!(-���,h��~���!��0|x[�s:�ǛC�w��7���IcVTZV����;{1��z$����n �A+W��v�w�(�>���`�/��_*N
���w�#��/�w�
��1} �e�Ns`W�Q\&h� �0~��:��ݳ`jo�K�#���m�-!!MH�N׃�6�V4�P��-�3	�W��z,Q�[���	�`wճ��ł���;�
o�+b����
O�|����(��##��:���(�W D���
Pt���9���������7ɲ7(���B��)Z�f�D����;��cWp�픈��B��ߛ�2~f����U�j=jf����cI�@���X���R����[������;���V��Bl��0�'�1�B�0LSMIΨ"�+;�p�/�E�LC��!A�{J	^�׎�yG;(�g�J��ƷM���̖�mԘ�k�a"˪J/qJq<�A�B��'�.�A&u�/��,��1-P@��5�`"�-"Ca��P�"#��2�7��-��)h�z���Y�Hsۈ0b:��l`�O�n�CX3