XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���n,A�*J�!��=ٯ�rb��Le���r�z�1�7�*��3�!���Ԟ�=f�/(5Ms��2歑�zX����K���M%���7�_��a���w��Mru�6��l���e"=�K(+ΰ�M9�5���ӭc�y��k��T4���uYځ��9�ǹ;�����68BTP������%"��>�Ƥ�l,���U�%+����ф%��c����Rn�-���ܧo���U��*�ڍ9�#8�r �����N�Qle}�j��<���0�)�/c�z@���u~=��P��n�&ԇnf�pJ��k��@���{>�z�����C�!r
Q4�k,��B�VfByr��/���؂U	�6�$QC�r�_uS�&\�;o
� �<݀�H-�#�1��bx�q����t��_���{DgZ���!Q�l*-6�[D<��4s�z��n�9ɚ����9`�Cr����]s�W���ϩ��@I�C�J��ٮ��B#�o��?��בgŅ���R�Q��r��$�p�F�����\-�N�wV_��|�?w�� �|@����i��x����I1g�K���	{h��X娎���
4��@��m9���Qx��}XҐś��J�75�d��#������V�%�J�S�QLȹ� %:?n!NM�O�3g7��-�|Z��Q,�_����8��!q�B�67�Q&L�����q�{*)�"BnL��1�A�����4���#�^T}J8�����Hӫ/A�?�;����7j�oXlxVHYEB    55a7     e50�H:#�-��Q�`8Ԥ�;��U�O>״w2�=�l1��a�S��SX��h��1Q�'�a!j5����ΰq��nޗ�<����"3�Y�Hm��	w�g�g-��<�y��J�`'����X��Pyw2�Hi�{`R�ʠ�H|\k�`N͛�� �djP���6,�-M)n����MB]q��h��-�L�QY#N��
5He\3aVv&{|'���̣lWb3�0���g�u�l�\����[(��`ݖ��1j���z��8~�Ƭ�qW��z�������κ�yF ���k� �y�G9�Z�+���ޜ;�^wj.���
sz�g��Oͧ�gg�"���e��lޝh&�C�2��h"�`�wT*Rw��b\��3uBz��{S�8c��p/�L���S_*��W�@�������qA�]�D�t��V�R9�L,�&��/4�ѯ��́�o�W������)CЉ���{:V�M�m���o~��:�+K�_,��L�[<����I�eH�D9?L7���kF;g��~.�19�l������9|��w��m ܾ2Uܼ2����H=�0����E������\���L�,K�
B��l���dN^��BZ�����ݞ(3mk�9\�T��p:H��O���q<��11�8�G���������΁_��U��� �/)�/AL	�TKܴ^� ��ҁ���N��s�Ll ��N)$�X��Q�4ofn}[x�o��#	E�[�@���t��%�kP��A�e@�T:��Z�}F� a��u���2n�?/o1��.ݎ�
7\��u{�g�1
,~QSdo����Tz[ߥ�(?}~ nj&Y|����k�2��J&��nh7{���987S��L�i{
��чEޗ�m����U�5��C���]�^>G���pt��:@ӂ�+�\]0-H�_6��%A���J�ԗ	��j���u�[ѥ��j�nE��`+DrtR#�zC�h炅�{h���9��C̅��9�_���F �j��&���pb1�y'Zk�ۯv)R:{��6AH�C���?ƽ��Fo� @�^I7���OK�@{�h ����~su�(�[9���&̨���T��g�~e-#Cw	�߶F�m�s�Z��xǄ1l� ��S{q��[��z\��3q���-^��xςg�O��	�na���{ln�8ܟB:M�N�)�X;��ke���b`j�Ć}'y��CK�����4T/JO?o`Sv��)׾!!��F��Ƚ�d^9�Ch !t6���/���+q��'F�J�i�?Q�m�i�������XQ#m�r޹���$���@�5���j}�銑@e��:>����@�>8�5��=(�2��H[Ձ�"�z���7s�!4G��/��������(�H첈j���W�Z��me���. ���3�Jŝ
K,р^�ſ�d-�yB���WL����	�)	y��TA����%ʝ�[߯@~��`��40X���{�R�G1�/^�b|jG_�7�/�ܯ���Ïn��Sڐ�*Ȫ�,c��
>�
r���i�v 
`�/ہ�=�J0,^�F�Sl�d#�M��r�\�<�"4�fAs�(�&�C�[�2ȍ���K9�w��O���wW�M�[�(�N�����^��N�\\Y=���U�n�AD!S¨Gz��[�Q�	UL|-������ԯ���`	V�A�����v%�hF�Z-��sNb�����f���{
`,YG�@$tK�<q�_$49%ytb����}��}/���3��o��C=/�o��ݏ>3�Զ��ĵH����[���wY�t����Z��{�Ab��
�2<AP����nƣ���������Lc����pC%�\�����Ao�]C�T� �;�֒��$���!��-���8�|��#�	:�`O˒����}��&�ʰ���K� �Y/��6녌k<��`S����^{/��D�|��5�/X��n�)dq�}����$kO#�RY`�����>�x�f&�L˪� T������];n�s�ؠ�F;l{�<ڥӉʥ�P5��RJ)~@$�E��I�8ev�;-�wq��
�#[�xu��@�Kq��Gd�=���d��d���PK���/�i`!��\�\��`!�?������u�Ņz���ZE^k� ����	׽.6g��'���(��17��݄Z)DZ|��V�M����t��w���^V�iih�2x̝�䄣N绍���*�:�hY�fB ��S�yo���8�Ц��_����A���@�?�d�j��heD�0�4�V+�;u�I�Y�.<��)%��f3��;O����j �{��S���F���$��������]��Z^Z֬>��(�zIJ �:[�[q�D�u�գ�Ru�`���q����j��,���:N{^��E��˪�&�M��36qA)H��f�4%J�]�� +P���X���>�P:p���G��&�	�0�+��r�청�.���^�����z�L�4���K8��L�ae�	�)�i��*�JNL*v��.�Yxq��)T� n/a�0�w݆P���`�j�]:�+/~œ�@����H��F���]
�O0�;ބ�w�HE�m���}��dY��Xc���ZM��yݙj�����J�nO��'�Fj�Ԣ��{��?��)P踏��tS%�B��E�cr(@�c;+רIht �_R5�\��zth���Kl�|�mT��2������ߵ���@猿{���x��&�y�_�x& ����ˣ�Ay;�O�J�[��q���(VV:�����*��f ���5R�F�;�,�y�����~�����W�AXI��D&��^����:A�1+C�UU��L܌n����y�B/�FliR����|l��`/X��������n�2	�K�%�Z/m�'����*�4��W�V�9d6��j��Z[q�Κ�a�wc*�s�n�U �	(2e�w�tM_��M<r�N�#�w�B���o���"���Ѐ�����8?����i�W)��J��ɷo�^݂��\rS�8=+(ju�9/3��'O#~��q;駗g8�T�M�i'���E����Fˢkp�}Y��{g��m$�KˢZw�Z�r�_@�9K)���*�"�K������dbp�=>,��Q����F��7E�?��f�-���<؞�����������Ι�Ca��R���A�c�)����/z#��p�31�)|:R�sU:�^�$������������3h��/���yJΤ}�w�sk��+v+�G)rNcD��I�r�Q��~�ۭf��f����dT�$U��??$���23Et�����q�C*�Z����Y�Iu}LU���?R�n��dE��V�l�%ݵ{���S4�W_��Lt�b.TVh�tUK���F)q�Y�;A�(��C6�۽@��R�
�A(9�J=�^z﹐vx()ܲ�K�
@�������n���r6�8es��d�L�K����6up�!Mm�J�C�Mˀ�ïi�(���}���[��,2we�F�w��PnB���
����;;�WfD��8��1p�]4C$N'���o������P�%��R� �d��*��Br��/d�}i��